----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date:     
-- Design Name: 
-- Module Name:     
-- Project Name: 
-- Target Devices: 
-- Tool versions: 
-- Description: 
--
-- Dependencies: 
--
-- Revision: 
-- Revision 0.01 - File Created
-- Additional Comments: 
--
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity TPG is
  Port (
    -- from clock wizard
    clk_in_100        : in  STD_LOGIC;
    clk_in_50         : in  STD_LOGIC;
    locked_in         : in  STD_LOGIC;
    -------------------------------------------------------
    test_data         : in  STD_LOGIC_VECTOR(11 downto 0);
    rom_adr           : out STD_LOGIC_VECTOR(16 downto 0);
    rom_dat           : in  STD_LOGIC_VECTOR(15 downto 0);
    -------------------------------------------------------
    mode_sel          : in STD_LOGIC_VECTOR( 3 downto 0);
    --vid interface to AXI-Stream @ 25MHz
    vid_data          : out std_logic_vector(23 downto 0);  -- RRRRRRRR BBBBBBBB GGGGGGGG
    vid_active_video  : out std_logic;
    vid_field_id      : out std_logic;
    vid_hsync         : out std_logic;
    vid_vsync         : out std_logic;
    -- zybo VGA interface 640x480 @ 25MHz
    RGB_data          : out STD_LOGIC_VECTOR(23 downto 0);
    Hsync             : out STD_LOGIC;
    Vsync             : out STD_LOGIC
  );
end TPG;


library UNISIM;
use UNISIM.VComponents.all;

architecture Structure of TPG is
  signal OVtpg_inst_VSYNC_60 : STD_LOGIC; 
  signal OVtpg_inst_HREF_61 : STD_LOGIC; 
  signal NlwRenamedSignal_SIF_inst_RGB_data_23_Q : STD_LOGIC; 
  signal NlwRenamedSignal_SIF_inst_RGB_data_22_Q : STD_LOGIC; 
  signal NlwRenamedSignal_SIF_inst_RGB_data_21_Q : STD_LOGIC; 
  signal NlwRenamedSignal_SIF_inst_RGB_data_20_Q : STD_LOGIC; 
  signal NlwRenamedSignal_SIF_inst_RGB_data_16_Q : STD_LOGIC; 
  signal NlwRenamedSignal_SIF_inst_RGB_data_15_Q : STD_LOGIC; 
  signal NlwRenamedSignal_SIF_inst_RGB_data_14_Q : STD_LOGIC; 
  signal NlwRenamedSignal_SIF_inst_RGB_data_13_Q : STD_LOGIC; 
  signal NlwRenamedSignal_SIF_inst_RGB_data_12_Q : STD_LOGIC; 
  signal NlwRenamedSignal_SIF_inst_RGB_data_11_Q : STD_LOGIC; 
  signal NlwRenamedSignal_SIF_inst_RGB_data_8_Q : STD_LOGIC; 
  signal NlwRenamedSignal_SIF_inst_RGB_data_7_Q : STD_LOGIC; 
  signal NlwRenamedSignal_SIF_inst_RGB_data_6_Q : STD_LOGIC; 
  signal NlwRenamedSignal_SIF_inst_RGB_data_5_Q : STD_LOGIC; 
  signal NlwRenamedSignal_SIF_inst_RGB_data_4_Q : STD_LOGIC; 
  signal NlwRenamedSignal_SIF_inst_RGB_data_0_Q : STD_LOGIC; 
  signal NlwRenamedSig_OI_SIF_inst_vid_active_video : STD_LOGIC; 
  signal NlwRenamedSig_OI_SIF_inst_Hsync : STD_LOGIC; 
  signal NlwRenamedSig_OI_SIF_inst_Vsync : STD_LOGIC; 
  signal MRST : STD_LOGIC; 
  signal NlwRenamedSig_OI_vid_field_id : STD_LOGIC; 
  signal N1 : STD_LOGIC; 
  signal OVtpg_inst_Mmux_pixel_out_12_pixel_out_23_mux_50_OUT3113 : STD_LOGIC; 
  signal OVtpg_inst_Mmux_pixel_out_12_pixel_out_23_mux_50_OUT3112 : STD_LOGIC; 
  signal OVtpg_inst_Mmux_pixel_out_12_pixel_out_23_mux_50_OUT3142 : STD_LOGIC; 
  signal OVtpg_inst_Mmux_pixel_out_12_pixel_out_23_mux_50_OUT4112 : STD_LOGIC; 
  signal OVtpg_inst_Mmux_pixel_out_12_pixel_out_23_mux_50_OUT3111 : STD_LOGIC; 
  signal OVtpg_inst_n02371 : STD_LOGIC; 
  signal OVtpg_inst_Col_10_GND_7_o_equal_4_o_10_1 : STD_LOGIC; 
  signal OVtpg_inst_Mmux_pixel_out_12_pixel_out_23_mux_50_OUT317 : STD_LOGIC; 
  signal OVtpg_inst_Mmux_pixel_out_12_pixel_out_23_mux_50_OUT15 : STD_LOGIC; 
  signal OVtpg_inst_Row_10_GND_7_o_equal_8_o_10_1 : STD_LOGIC; 
  signal OVtpg_inst_Row_10_GND_7_o_equal_5_o_10_1_96 : STD_LOGIC; 
  signal OVtpg_inst_n0315_inv1 : STD_LOGIC; 
  signal OVtpg_inst_Mmux_pixel_out_12_pixel_out_23_mux_50_OUT316 : STD_LOGIC; 
  signal OVtpg_inst_Result_10_2 : STD_LOGIC; 
  signal OVtpg_inst_Result_9_2 : STD_LOGIC; 
  signal OVtpg_inst_Result_8_2 : STD_LOGIC; 
  signal OVtpg_inst_Result_7_2 : STD_LOGIC; 
  signal OVtpg_inst_Result_6_2 : STD_LOGIC; 
  signal OVtpg_inst_Result_5_2 : STD_LOGIC; 
  signal OVtpg_inst_Result_4_2 : STD_LOGIC; 
  signal OVtpg_inst_Result_3_2 : STD_LOGIC; 
  signal OVtpg_inst_Result_2_2 : STD_LOGIC; 
  signal OVtpg_inst_Result_1_3 : STD_LOGIC; 
  signal OVtpg_inst_Result_0_3 : STD_LOGIC; 
  signal OVtpg_inst_Mcount_Col_val : STD_LOGIC; 
  signal OVtpg_inst_Result_10_1 : STD_LOGIC; 
  signal OVtpg_inst_Result_9_1 : STD_LOGIC; 
  signal OVtpg_inst_Result_8_1 : STD_LOGIC; 
  signal OVtpg_inst_Result_7_1 : STD_LOGIC; 
  signal OVtpg_inst_Result_6_1 : STD_LOGIC; 
  signal OVtpg_inst_Result_5_1 : STD_LOGIC; 
  signal OVtpg_inst_Result_4_1 : STD_LOGIC; 
  signal OVtpg_inst_Result_3_1 : STD_LOGIC; 
  signal OVtpg_inst_Result_2_1 : STD_LOGIC; 
  signal OVtpg_inst_Result_1_2 : STD_LOGIC; 
  signal OVtpg_inst_Result_0_2 : STD_LOGIC; 
  signal OVtpg_inst_Mcount_Row_val : STD_LOGIC; 
  signal OVtpg_inst_Result_1_1 : STD_LOGIC; 
  signal OVtpg_inst_Result_0_1 : STD_LOGIC; 
  signal OVtpg_inst_n0395_inv : STD_LOGIC; 
  signal OVtpg_inst_Mram_MODE_3_PWR_7_o_wide_mux_9_OUT2 : STD_LOGIC; 
  signal OVtpg_inst_Mram_MODE_3_PWR_7_o_wide_mux_9_OUT1 : STD_LOGIC; 
  signal OVtpg_inst_Mram_MODE_3_PWR_7_o_wide_mux_9_OUT : STD_LOGIC; 
  signal OVtpg_inst_n0358_inv_184 : STD_LOGIC; 
  signal OVtpg_inst_pixel_out_12_pixel_out_23_mux_50_OUT_0_Q : STD_LOGIC; 
  signal OVtpg_inst_pixel_out_12_pixel_out_23_mux_50_OUT_1_Q : STD_LOGIC; 
  signal OVtpg_inst_pixel_out_12_pixel_out_23_mux_50_OUT_2_Q : STD_LOGIC; 
  signal OVtpg_inst_pixel_out_12_pixel_out_23_mux_50_OUT_3_Q : STD_LOGIC; 
  signal OVtpg_inst_pixel_out_12_pixel_out_23_mux_50_OUT_4_Q : STD_LOGIC; 
  signal OVtpg_inst_pixel_out_12_pixel_out_23_mux_50_OUT_5_Q : STD_LOGIC; 
  signal OVtpg_inst_pixel_out_12_pixel_out_23_mux_50_OUT_6_Q : STD_LOGIC; 
  signal OVtpg_inst_pixel_out_12_pixel_out_23_mux_50_OUT_7_Q : STD_LOGIC; 
  signal OVtpg_inst_Col_10_GND_7_o_equal_4_o : STD_LOGIC; 
  signal OVtpg_inst_Inside : STD_LOGIC; 
  signal OVtpg_inst_n0270 : STD_LOGIC; 
  signal OVtpg_inst_Cen : STD_LOGIC; 
  signal OVtpg_inst_PCLK : STD_LOGIC; 
  signal OVtpg_inst_n0244_198 : STD_LOGIC; 
  signal OVtpg_inst_n0254_199 : STD_LOGIC; 
  signal OVtpg_inst_n0262_200 : STD_LOGIC; 
  signal OVtpg_inst_Hsynci_234 : STD_LOGIC; 
  signal OVtpg_inst_Active_235 : STD_LOGIC; 
  signal OVtpg_inst_Hrefi_236 : STD_LOGIC; 
  signal OVtpg_inst_Vsynci_237 : STD_LOGIC; 
  signal OVtpg_inst_Row_10_PWR_7_o_div_45_o_0_12 : STD_LOGIC; 
  signal OVtpg_inst_Row_10_PWR_7_o_div_45_o_0_11 : STD_LOGIC; 
  signal OVtpg_inst_Row_10_PWR_7_o_div_45_Madd_a_10_GND_9_o_add_19_OUT_10_0_lut_7_Q : STD_LOGIC; 
  signal OVtpg_inst_Row_10_PWR_7_o_div_45_Madd_a_10_GND_9_o_add_19_OUT_10_0_lut_6_Q : STD_LOGIC; 
  signal OVtpg_inst_Row_10_PWR_7_o_div_45_n0441_8_Q : STD_LOGIC; 
  signal OVtpg_inst_Col_10_PWR_7_o_div_44_o_0_13 : STD_LOGIC; 
  signal OVtpg_inst_Col_10_PWR_7_o_div_44_Madd_a_10_GND_8_o_add_21_OUT_10_0_lut_7_Q : STD_LOGIC; 
  signal SIF_inst_Reset_OR_DriverANDClockEnable : STD_LOGIC; 
  signal SIF_inst_oddpix1 : STD_LOGIC; 
  signal SIF_inst_n0060_inv : STD_LOGIC; 
  signal SIF_inst_oddpix_INV_358_o : STD_LOGIC; 
  signal SIF_inst_VS_in_INV_360_o : STD_LOGIC; 
  signal SIF_inst_oddpix_252 : STD_LOGIC; 
  signal OVtpg_inst_Mmux_pixel_out_12_pixel_out_23_mux_50_OUT3171_261 : STD_LOGIC; 
  signal OVtpg_inst_Mmux_pixel_out_12_pixel_out_23_mux_50_OUT3172_262 : STD_LOGIC; 
  signal OVtpg_inst_Mmux_pixel_out_12_pixel_out_23_mux_50_OUT3173_263 : STD_LOGIC; 
  signal OVtpg_inst_Mmux_pixel_out_12_pixel_out_23_mux_50_OUT3177_264 : STD_LOGIC; 
  signal OVtpg_inst_Mmux_pixel_out_12_pixel_out_23_mux_50_OUT3178_265 : STD_LOGIC; 
  signal OVtpg_inst_Mmux_pixel_out_12_pixel_out_23_mux_50_OUT41121_266 : STD_LOGIC; 
  signal OVtpg_inst_Mmux_pixel_out_12_pixel_out_23_mux_50_OUT41122_267 : STD_LOGIC; 
  signal OVtpg_inst_Mmux_pixel_out_12_pixel_out_23_mux_50_OUT41123_268 : STD_LOGIC; 
  signal OVtpg_inst_Mmux_pixel_out_12_pixel_out_23_mux_50_OUT41124_269 : STD_LOGIC; 
  signal OVtpg_inst_Mmux_pixel_out_12_pixel_out_23_mux_50_OUT41126_270 : STD_LOGIC; 
  signal OVtpg_inst_Mmux_pixel_out_12_pixel_out_23_mux_50_OUT41128_271 : STD_LOGIC; 
  signal N4 : STD_LOGIC; 
  signal N6 : STD_LOGIC; 
  signal N8 : STD_LOGIC; 
  signal OVtpg_inst_n0395_inv3_275 : STD_LOGIC; 
  signal OVtpg_inst_Mmux_pixel_out_12_pixel_out_23_mux_50_OUT7 : STD_LOGIC; 
  signal OVtpg_inst_Mmux_pixel_out_12_pixel_out_23_mux_50_OUT71_277 : STD_LOGIC; 
  signal OVtpg_inst_Mmux_pixel_out_12_pixel_out_23_mux_50_OUT6 : STD_LOGIC; 
  signal OVtpg_inst_Mmux_pixel_out_12_pixel_out_23_mux_50_OUT61_279 : STD_LOGIC; 
  signal OVtpg_inst_Mmux_pixel_out_12_pixel_out_23_mux_50_OUT8 : STD_LOGIC; 
  signal N10 : STD_LOGIC; 
  signal N12 : STD_LOGIC; 
  signal N14 : STD_LOGIC; 
  signal N16 : STD_LOGIC; 
  signal OVtpg_inst_Mmux_pixel_out_12_pixel_out_23_mux_50_OUT3 : STD_LOGIC; 
  signal OVtpg_inst_Mmux_pixel_out_12_pixel_out_23_mux_50_OUT31_286 : STD_LOGIC; 
  signal OVtpg_inst_Inside1_287 : STD_LOGIC; 
  signal OVtpg_inst_Inside2_288 : STD_LOGIC; 
  signal N18 : STD_LOGIC; 
  signal N20 : STD_LOGIC; 
  signal OVtpg_inst_Mmux_pixel_out_12_pixel_out_23_mux_50_OUT3161_291 : STD_LOGIC; 
  signal OVtpg_inst_Mmux_pixel_out_12_pixel_out_23_mux_50_OUT3162_292 : STD_LOGIC; 
  signal OVtpg_inst_Mmux_pixel_out_12_pixel_out_23_mux_50_OUT3163_293 : STD_LOGIC; 
  signal OVtpg_inst_Mmux_pixel_out_12_pixel_out_23_mux_50_OUT3164 : STD_LOGIC; 
  signal OVtpg_inst_Mmux_pixel_out_12_pixel_out_23_mux_50_OUT3165_295 : STD_LOGIC; 
  signal OVtpg_inst_Mmux_pixel_out_12_pixel_out_23_mux_50_OUT3166_296 : STD_LOGIC; 
  signal OVtpg_inst_Mmux_pixel_out_12_pixel_out_23_mux_50_OUT3167_297 : STD_LOGIC; 
  signal OVtpg_inst_Mmux_pixel_out_12_pixel_out_23_mux_50_OUT3169_298 : STD_LOGIC; 
  signal OVtpg_inst_Hsynci_glue_set_299 : STD_LOGIC; 
  signal OVtpg_inst_Active_glue_set_300 : STD_LOGIC; 
  signal OVtpg_inst_Hrefi_glue_set_301 : STD_LOGIC; 
  signal OVtpg_inst_Vsynci_glue_set : STD_LOGIC; 
  signal SIF_inst_vid_active_video_glue_set_303 : STD_LOGIC; 
  signal OVtpg_inst_Mcount_Col_cy_9_rt_304 : STD_LOGIC; 
  signal OVtpg_inst_Mcount_Col_cy_8_rt_305 : STD_LOGIC; 
  signal OVtpg_inst_Mcount_Col_cy_7_rt_306 : STD_LOGIC; 
  signal OVtpg_inst_Mcount_Col_cy_6_rt_307 : STD_LOGIC; 
  signal OVtpg_inst_Mcount_Col_cy_5_rt_308 : STD_LOGIC; 
  signal OVtpg_inst_Mcount_Col_cy_4_rt_309 : STD_LOGIC; 
  signal OVtpg_inst_Mcount_Col_cy_3_rt_310 : STD_LOGIC; 
  signal OVtpg_inst_Mcount_Col_cy_2_rt_311 : STD_LOGIC; 
  signal OVtpg_inst_Mcount_Col_cy_1_rt_312 : STD_LOGIC; 
  signal OVtpg_inst_Mcount_Row_cy_9_rt_313 : STD_LOGIC; 
  signal OVtpg_inst_Mcount_Row_cy_8_rt_314 : STD_LOGIC; 
  signal OVtpg_inst_Mcount_Row_cy_7_rt_315 : STD_LOGIC; 
  signal OVtpg_inst_Mcount_Row_cy_6_rt_316 : STD_LOGIC; 
  signal OVtpg_inst_Mcount_Row_cy_5_rt_317 : STD_LOGIC; 
  signal OVtpg_inst_Mcount_Row_cy_4_rt_318 : STD_LOGIC; 
  signal OVtpg_inst_Mcount_Row_cy_3_rt_319 : STD_LOGIC; 
  signal OVtpg_inst_Mcount_Row_cy_2_rt_320 : STD_LOGIC; 
  signal OVtpg_inst_Mcount_Row_cy_1_rt_321 : STD_LOGIC; 
  signal OVtpg_inst_Mcount_addr_cy_15_rt_322 : STD_LOGIC; 
  signal OVtpg_inst_Mcount_addr_cy_14_rt_323 : STD_LOGIC; 
  signal OVtpg_inst_Mcount_addr_cy_13_rt_324 : STD_LOGIC; 
  signal OVtpg_inst_Mcount_addr_cy_12_rt_325 : STD_LOGIC; 
  signal OVtpg_inst_Mcount_addr_cy_11_rt_326 : STD_LOGIC; 
  signal OVtpg_inst_Mcount_addr_cy_10_rt_327 : STD_LOGIC; 
  signal OVtpg_inst_Mcount_addr_cy_9_rt_328 : STD_LOGIC; 
  signal OVtpg_inst_Mcount_addr_cy_8_rt_329 : STD_LOGIC; 
  signal OVtpg_inst_Mcount_addr_cy_7_rt_330 : STD_LOGIC; 
  signal OVtpg_inst_Mcount_addr_cy_6_rt_331 : STD_LOGIC; 
  signal OVtpg_inst_Mcount_addr_cy_5_rt_332 : STD_LOGIC; 
  signal OVtpg_inst_Mcount_addr_cy_4_rt_333 : STD_LOGIC; 
  signal OVtpg_inst_Mcount_addr_cy_3_rt_334 : STD_LOGIC; 
  signal OVtpg_inst_Mcount_addr_cy_2_rt_335 : STD_LOGIC; 
  signal OVtpg_inst_Mcount_addr_cy_1_rt_336 : STD_LOGIC; 
  signal OVtpg_inst_Mcount_Col_xor_10_rt_337 : STD_LOGIC; 
  signal OVtpg_inst_Mcount_Row_xor_10_rt_338 : STD_LOGIC; 
  signal N22 : STD_LOGIC; 
  signal N32 : STD_LOGIC; 
  signal N33 : STD_LOGIC; 
  signal N35 : STD_LOGIC; 
  signal N36 : STD_LOGIC; 
  signal N39 : STD_LOGIC; 
  signal N42 : STD_LOGIC; 
  signal N44 : STD_LOGIC; 
  signal N48 : STD_LOGIC; 
  signal N49 : STD_LOGIC; 
  signal N55 : STD_LOGIC; 
  signal N56 : STD_LOGIC; 
  signal N91 : STD_LOGIC; 
  signal N92 : STD_LOGIC; 
  signal N94 : STD_LOGIC; 
  signal N95 : STD_LOGIC; 
  signal N97 : STD_LOGIC; 
  signal N98 : STD_LOGIC; 
  signal N100 : STD_LOGIC; 
  signal N101 : STD_LOGIC; 
  signal N102 : STD_LOGIC; 
  signal N103 : STD_LOGIC; 
  signal N105 : STD_LOGIC; 
  signal N106 : STD_LOGIC; 
  signal N107 : STD_LOGIC; 
  signal N108 : STD_LOGIC; 
  signal N110 : STD_LOGIC; 
  signal N111 : STD_LOGIC; 
  signal N112 : STD_LOGIC; 
  signal N114 : STD_LOGIC; 
  signal N115 : STD_LOGIC; 
  signal N116 : STD_LOGIC; 
  signal N124 : STD_LOGIC; 
  signal N125 : STD_LOGIC; 
  signal N126 : STD_LOGIC; 
  signal N127 : STD_LOGIC; 
  signal N128 : STD_LOGIC; 
  signal N129 : STD_LOGIC; 
  signal N130 : STD_LOGIC; 
  signal N131 : STD_LOGIC; 
  signal N132 : STD_LOGIC; 
  signal N134 : STD_LOGIC; 
  signal N136 : STD_LOGIC; 
  signal N137 : STD_LOGIC; 
  signal N138 : STD_LOGIC; 
  signal N139 : STD_LOGIC; 
  signal N140 : STD_LOGIC; 
  signal N141 : STD_LOGIC; 
  signal N143 : STD_LOGIC; 
  signal NlwRenamedSig_OI_OVtpg_inst_addr : STD_LOGIC_VECTOR ( 16 downto 0 ); 
  signal OVtpg_inst_D : STD_LOGIC_VECTOR ( 7 downto 0 ); 
  signal OVtpg_inst_Mcount_Col_cy : STD_LOGIC_VECTOR ( 9 downto 0 ); 
  signal OVtpg_inst_Mcount_Col_lut : STD_LOGIC_VECTOR ( 0 downto 0 ); 
  signal OVtpg_inst_Mcount_Row_cy : STD_LOGIC_VECTOR ( 9 downto 0 ); 
  signal OVtpg_inst_Mcount_Row_lut : STD_LOGIC_VECTOR ( 0 downto 0 ); 
  signal OVtpg_inst_Mcount_addr_cy : STD_LOGIC_VECTOR ( 15 downto 0 ); 
  signal OVtpg_inst_Mcount_addr_lut : STD_LOGIC_VECTOR ( 0 downto 0 ); 
  signal OVtpg_inst_Result : STD_LOGIC_VECTOR ( 16 downto 1 ); 
  signal OVtpg_inst_n0133 : STD_LOGIC_VECTOR ( 3 downto 0 ); 
  signal OVtpg_inst_n0134 : STD_LOGIC_VECTOR ( 3 downto 0 ); 
  signal OVtpg_inst_Col : STD_LOGIC_VECTOR ( 10 downto 0 ); 
  signal OVtpg_inst_Row : STD_LOGIC_VECTOR ( 10 downto 0 ); 
  signal OVtpg_inst_pmode : STD_LOGIC_VECTOR ( 2 downto 0 ); 
  signal OVtpg_inst_ClkDiv : STD_LOGIC_VECTOR ( 1 downto 0 ); 
  signal SIF_inst_FirstByte : STD_LOGIC_VECTOR ( 7 downto 0 ); 
begin
  rom_adr(16) <= NlwRenamedSig_OI_OVtpg_inst_addr(16);
  rom_adr(15) <= NlwRenamedSig_OI_OVtpg_inst_addr(15);
  rom_adr(14) <= NlwRenamedSig_OI_OVtpg_inst_addr(14);
  rom_adr(13) <= NlwRenamedSig_OI_OVtpg_inst_addr(13);
  rom_adr(12) <= NlwRenamedSig_OI_OVtpg_inst_addr(12);
  rom_adr(11) <= NlwRenamedSig_OI_OVtpg_inst_addr(11);
  rom_adr(10) <= NlwRenamedSig_OI_OVtpg_inst_addr(10);
  rom_adr(9) <= NlwRenamedSig_OI_OVtpg_inst_addr(9);
  rom_adr(8) <= NlwRenamedSig_OI_OVtpg_inst_addr(8);
  rom_adr(7) <= NlwRenamedSig_OI_OVtpg_inst_addr(7);
  rom_adr(6) <= NlwRenamedSig_OI_OVtpg_inst_addr(6);
  rom_adr(5) <= NlwRenamedSig_OI_OVtpg_inst_addr(5);
  rom_adr(4) <= NlwRenamedSig_OI_OVtpg_inst_addr(4);
  rom_adr(3) <= NlwRenamedSig_OI_OVtpg_inst_addr(3);
  rom_adr(2) <= NlwRenamedSig_OI_OVtpg_inst_addr(2);
  rom_adr(1) <= NlwRenamedSig_OI_OVtpg_inst_addr(1);
  rom_adr(0) <= NlwRenamedSig_OI_OVtpg_inst_addr(0);
  vid_data(23) <= NlwRenamedSignal_SIF_inst_RGB_data_23_Q;
  vid_data(22) <= NlwRenamedSignal_SIF_inst_RGB_data_22_Q;
  vid_data(21) <= NlwRenamedSignal_SIF_inst_RGB_data_21_Q;
  vid_data(20) <= NlwRenamedSignal_SIF_inst_RGB_data_20_Q;
  vid_data(19) <= NlwRenamedSignal_SIF_inst_RGB_data_16_Q;
  vid_data(18) <= NlwRenamedSignal_SIF_inst_RGB_data_16_Q;
  vid_data(17) <= NlwRenamedSignal_SIF_inst_RGB_data_16_Q;
  vid_data(16) <= NlwRenamedSignal_SIF_inst_RGB_data_16_Q;
  vid_data(15) <= NlwRenamedSignal_SIF_inst_RGB_data_7_Q;
  vid_data(14) <= NlwRenamedSignal_SIF_inst_RGB_data_6_Q;
  vid_data(13) <= NlwRenamedSignal_SIF_inst_RGB_data_5_Q;
  vid_data(12) <= NlwRenamedSignal_SIF_inst_RGB_data_4_Q;
  vid_data(11) <= NlwRenamedSignal_SIF_inst_RGB_data_0_Q;
  vid_data(10) <= NlwRenamedSignal_SIF_inst_RGB_data_0_Q;
  vid_data(9) <= NlwRenamedSignal_SIF_inst_RGB_data_0_Q;
  vid_data(8) <= NlwRenamedSignal_SIF_inst_RGB_data_0_Q;
  vid_data(7) <= NlwRenamedSignal_SIF_inst_RGB_data_15_Q;
  vid_data(6) <= NlwRenamedSignal_SIF_inst_RGB_data_14_Q;
  vid_data(5) <= NlwRenamedSignal_SIF_inst_RGB_data_13_Q;
  vid_data(4) <= NlwRenamedSignal_SIF_inst_RGB_data_12_Q;
  vid_data(3) <= NlwRenamedSignal_SIF_inst_RGB_data_11_Q;
  vid_data(2) <= NlwRenamedSignal_SIF_inst_RGB_data_8_Q;
  vid_data(1) <= NlwRenamedSignal_SIF_inst_RGB_data_8_Q;
  vid_data(0) <= NlwRenamedSignal_SIF_inst_RGB_data_8_Q;
  RGB_data(23) <= NlwRenamedSignal_SIF_inst_RGB_data_23_Q;
  RGB_data(22) <= NlwRenamedSignal_SIF_inst_RGB_data_22_Q;
  RGB_data(21) <= NlwRenamedSignal_SIF_inst_RGB_data_21_Q;
  RGB_data(20) <= NlwRenamedSignal_SIF_inst_RGB_data_20_Q;
  RGB_data(19) <= NlwRenamedSignal_SIF_inst_RGB_data_16_Q;
  RGB_data(18) <= NlwRenamedSignal_SIF_inst_RGB_data_16_Q;
  RGB_data(17) <= NlwRenamedSignal_SIF_inst_RGB_data_16_Q;
  RGB_data(16) <= NlwRenamedSignal_SIF_inst_RGB_data_16_Q;
  RGB_data(15) <= NlwRenamedSignal_SIF_inst_RGB_data_15_Q;
  RGB_data(14) <= NlwRenamedSignal_SIF_inst_RGB_data_14_Q;
  RGB_data(13) <= NlwRenamedSignal_SIF_inst_RGB_data_13_Q;
  RGB_data(12) <= NlwRenamedSignal_SIF_inst_RGB_data_12_Q;
  RGB_data(11) <= NlwRenamedSignal_SIF_inst_RGB_data_11_Q;
  RGB_data(10) <= NlwRenamedSignal_SIF_inst_RGB_data_8_Q;
  RGB_data(9) <= NlwRenamedSignal_SIF_inst_RGB_data_8_Q;
  RGB_data(8) <= NlwRenamedSignal_SIF_inst_RGB_data_8_Q;
  RGB_data(7) <= NlwRenamedSignal_SIF_inst_RGB_data_7_Q;
  RGB_data(6) <= NlwRenamedSignal_SIF_inst_RGB_data_6_Q;
  RGB_data(5) <= NlwRenamedSignal_SIF_inst_RGB_data_5_Q;
  RGB_data(4) <= NlwRenamedSignal_SIF_inst_RGB_data_4_Q;
  RGB_data(3) <= NlwRenamedSignal_SIF_inst_RGB_data_0_Q;
  RGB_data(2) <= NlwRenamedSignal_SIF_inst_RGB_data_0_Q;
  RGB_data(1) <= NlwRenamedSignal_SIF_inst_RGB_data_0_Q;
  RGB_data(0) <= NlwRenamedSignal_SIF_inst_RGB_data_0_Q;
  vid_active_video <= NlwRenamedSig_OI_SIF_inst_vid_active_video;
  vid_field_id <= NlwRenamedSig_OI_vid_field_id;
  Hsync <= NlwRenamedSig_OI_SIF_inst_Hsync;
  Vsync <= NlwRenamedSig_OI_SIF_inst_Vsync;
  XST_GND : GND
    port map (
      G => NlwRenamedSig_OI_vid_field_id
    );
  XST_VCC : VCC
    port map (
      P => N1
    );
  OVtpg_inst_Mcount_Col_xor_10_Q : XORCY
    port map (
      CI => OVtpg_inst_Mcount_Col_cy(9),
      LI => OVtpg_inst_Mcount_Col_xor_10_rt_337,
      O => OVtpg_inst_Result_10_2
    );
  OVtpg_inst_Mcount_Col_xor_9_Q : XORCY
    port map (
      CI => OVtpg_inst_Mcount_Col_cy(8),
      LI => OVtpg_inst_Mcount_Col_cy_9_rt_304,
      O => OVtpg_inst_Result_9_2
    );
  OVtpg_inst_Mcount_Col_cy_9_Q : MUXCY
    port map (
      CI => OVtpg_inst_Mcount_Col_cy(8),
      DI => NlwRenamedSig_OI_vid_field_id,
      S => OVtpg_inst_Mcount_Col_cy_9_rt_304,
      O => OVtpg_inst_Mcount_Col_cy(9)
    );
  OVtpg_inst_Mcount_Col_xor_8_Q : XORCY
    port map (
      CI => OVtpg_inst_Mcount_Col_cy(7),
      LI => OVtpg_inst_Mcount_Col_cy_8_rt_305,
      O => OVtpg_inst_Result_8_2
    );
  OVtpg_inst_Mcount_Col_cy_8_Q : MUXCY
    port map (
      CI => OVtpg_inst_Mcount_Col_cy(7),
      DI => NlwRenamedSig_OI_vid_field_id,
      S => OVtpg_inst_Mcount_Col_cy_8_rt_305,
      O => OVtpg_inst_Mcount_Col_cy(8)
    );
  OVtpg_inst_Mcount_Col_xor_7_Q : XORCY
    port map (
      CI => OVtpg_inst_Mcount_Col_cy(6),
      LI => OVtpg_inst_Mcount_Col_cy_7_rt_306,
      O => OVtpg_inst_Result_7_2
    );
  OVtpg_inst_Mcount_Col_cy_7_Q : MUXCY
    port map (
      CI => OVtpg_inst_Mcount_Col_cy(6),
      DI => NlwRenamedSig_OI_vid_field_id,
      S => OVtpg_inst_Mcount_Col_cy_7_rt_306,
      O => OVtpg_inst_Mcount_Col_cy(7)
    );
  OVtpg_inst_Mcount_Col_xor_6_Q : XORCY
    port map (
      CI => OVtpg_inst_Mcount_Col_cy(5),
      LI => OVtpg_inst_Mcount_Col_cy_6_rt_307,
      O => OVtpg_inst_Result_6_2
    );
  OVtpg_inst_Mcount_Col_cy_6_Q : MUXCY
    port map (
      CI => OVtpg_inst_Mcount_Col_cy(5),
      DI => NlwRenamedSig_OI_vid_field_id,
      S => OVtpg_inst_Mcount_Col_cy_6_rt_307,
      O => OVtpg_inst_Mcount_Col_cy(6)
    );
  OVtpg_inst_Mcount_Col_xor_5_Q : XORCY
    port map (
      CI => OVtpg_inst_Mcount_Col_cy(4),
      LI => OVtpg_inst_Mcount_Col_cy_5_rt_308,
      O => OVtpg_inst_Result_5_2
    );
  OVtpg_inst_Mcount_Col_cy_5_Q : MUXCY
    port map (
      CI => OVtpg_inst_Mcount_Col_cy(4),
      DI => NlwRenamedSig_OI_vid_field_id,
      S => OVtpg_inst_Mcount_Col_cy_5_rt_308,
      O => OVtpg_inst_Mcount_Col_cy(5)
    );
  OVtpg_inst_Mcount_Col_xor_4_Q : XORCY
    port map (
      CI => OVtpg_inst_Mcount_Col_cy(3),
      LI => OVtpg_inst_Mcount_Col_cy_4_rt_309,
      O => OVtpg_inst_Result_4_2
    );
  OVtpg_inst_Mcount_Col_cy_4_Q : MUXCY
    port map (
      CI => OVtpg_inst_Mcount_Col_cy(3),
      DI => NlwRenamedSig_OI_vid_field_id,
      S => OVtpg_inst_Mcount_Col_cy_4_rt_309,
      O => OVtpg_inst_Mcount_Col_cy(4)
    );
  OVtpg_inst_Mcount_Col_xor_3_Q : XORCY
    port map (
      CI => OVtpg_inst_Mcount_Col_cy(2),
      LI => OVtpg_inst_Mcount_Col_cy_3_rt_310,
      O => OVtpg_inst_Result_3_2
    );
  OVtpg_inst_Mcount_Col_cy_3_Q : MUXCY
    port map (
      CI => OVtpg_inst_Mcount_Col_cy(2),
      DI => NlwRenamedSig_OI_vid_field_id,
      S => OVtpg_inst_Mcount_Col_cy_3_rt_310,
      O => OVtpg_inst_Mcount_Col_cy(3)
    );
  OVtpg_inst_Mcount_Col_xor_2_Q : XORCY
    port map (
      CI => OVtpg_inst_Mcount_Col_cy(1),
      LI => OVtpg_inst_Mcount_Col_cy_2_rt_311,
      O => OVtpg_inst_Result_2_2
    );
  OVtpg_inst_Mcount_Col_cy_2_Q : MUXCY
    port map (
      CI => OVtpg_inst_Mcount_Col_cy(1),
      DI => NlwRenamedSig_OI_vid_field_id,
      S => OVtpg_inst_Mcount_Col_cy_2_rt_311,
      O => OVtpg_inst_Mcount_Col_cy(2)
    );
  OVtpg_inst_Mcount_Col_xor_1_Q : XORCY
    port map (
      CI => OVtpg_inst_Mcount_Col_cy(0),
      LI => OVtpg_inst_Mcount_Col_cy_1_rt_312,
      O => OVtpg_inst_Result_1_3
    );
  OVtpg_inst_Mcount_Col_cy_1_Q : MUXCY
    port map (
      CI => OVtpg_inst_Mcount_Col_cy(0),
      DI => NlwRenamedSig_OI_vid_field_id,
      S => OVtpg_inst_Mcount_Col_cy_1_rt_312,
      O => OVtpg_inst_Mcount_Col_cy(1)
    );
  OVtpg_inst_Mcount_Col_xor_0_Q : XORCY
    port map (
      CI => NlwRenamedSig_OI_vid_field_id,
      LI => OVtpg_inst_Mcount_Col_lut(0),
      O => OVtpg_inst_Result_0_3
    );
  OVtpg_inst_Mcount_Col_cy_0_Q : MUXCY
    port map (
      CI => NlwRenamedSig_OI_vid_field_id,
      DI => N1,
      S => OVtpg_inst_Mcount_Col_lut(0),
      O => OVtpg_inst_Mcount_Col_cy(0)
    );
  OVtpg_inst_Mcount_Row_xor_10_Q : XORCY
    port map (
      CI => OVtpg_inst_Mcount_Row_cy(9),
      LI => OVtpg_inst_Mcount_Row_xor_10_rt_338,
      O => OVtpg_inst_Result_10_1
    );
  OVtpg_inst_Mcount_Row_xor_9_Q : XORCY
    port map (
      CI => OVtpg_inst_Mcount_Row_cy(8),
      LI => OVtpg_inst_Mcount_Row_cy_9_rt_313,
      O => OVtpg_inst_Result_9_1
    );
  OVtpg_inst_Mcount_Row_cy_9_Q : MUXCY
    port map (
      CI => OVtpg_inst_Mcount_Row_cy(8),
      DI => NlwRenamedSig_OI_vid_field_id,
      S => OVtpg_inst_Mcount_Row_cy_9_rt_313,
      O => OVtpg_inst_Mcount_Row_cy(9)
    );
  OVtpg_inst_Mcount_Row_xor_8_Q : XORCY
    port map (
      CI => OVtpg_inst_Mcount_Row_cy(7),
      LI => OVtpg_inst_Mcount_Row_cy_8_rt_314,
      O => OVtpg_inst_Result_8_1
    );
  OVtpg_inst_Mcount_Row_cy_8_Q : MUXCY
    port map (
      CI => OVtpg_inst_Mcount_Row_cy(7),
      DI => NlwRenamedSig_OI_vid_field_id,
      S => OVtpg_inst_Mcount_Row_cy_8_rt_314,
      O => OVtpg_inst_Mcount_Row_cy(8)
    );
  OVtpg_inst_Mcount_Row_xor_7_Q : XORCY
    port map (
      CI => OVtpg_inst_Mcount_Row_cy(6),
      LI => OVtpg_inst_Mcount_Row_cy_7_rt_315,
      O => OVtpg_inst_Result_7_1
    );
  OVtpg_inst_Mcount_Row_cy_7_Q : MUXCY
    port map (
      CI => OVtpg_inst_Mcount_Row_cy(6),
      DI => NlwRenamedSig_OI_vid_field_id,
      S => OVtpg_inst_Mcount_Row_cy_7_rt_315,
      O => OVtpg_inst_Mcount_Row_cy(7)
    );
  OVtpg_inst_Mcount_Row_xor_6_Q : XORCY
    port map (
      CI => OVtpg_inst_Mcount_Row_cy(5),
      LI => OVtpg_inst_Mcount_Row_cy_6_rt_316,
      O => OVtpg_inst_Result_6_1
    );
  OVtpg_inst_Mcount_Row_cy_6_Q : MUXCY
    port map (
      CI => OVtpg_inst_Mcount_Row_cy(5),
      DI => NlwRenamedSig_OI_vid_field_id,
      S => OVtpg_inst_Mcount_Row_cy_6_rt_316,
      O => OVtpg_inst_Mcount_Row_cy(6)
    );
  OVtpg_inst_Mcount_Row_xor_5_Q : XORCY
    port map (
      CI => OVtpg_inst_Mcount_Row_cy(4),
      LI => OVtpg_inst_Mcount_Row_cy_5_rt_317,
      O => OVtpg_inst_Result_5_1
    );
  OVtpg_inst_Mcount_Row_cy_5_Q : MUXCY
    port map (
      CI => OVtpg_inst_Mcount_Row_cy(4),
      DI => NlwRenamedSig_OI_vid_field_id,
      S => OVtpg_inst_Mcount_Row_cy_5_rt_317,
      O => OVtpg_inst_Mcount_Row_cy(5)
    );
  OVtpg_inst_Mcount_Row_xor_4_Q : XORCY
    port map (
      CI => OVtpg_inst_Mcount_Row_cy(3),
      LI => OVtpg_inst_Mcount_Row_cy_4_rt_318,
      O => OVtpg_inst_Result_4_1
    );
  OVtpg_inst_Mcount_Row_cy_4_Q : MUXCY
    port map (
      CI => OVtpg_inst_Mcount_Row_cy(3),
      DI => NlwRenamedSig_OI_vid_field_id,
      S => OVtpg_inst_Mcount_Row_cy_4_rt_318,
      O => OVtpg_inst_Mcount_Row_cy(4)
    );
  OVtpg_inst_Mcount_Row_xor_3_Q : XORCY
    port map (
      CI => OVtpg_inst_Mcount_Row_cy(2),
      LI => OVtpg_inst_Mcount_Row_cy_3_rt_319,
      O => OVtpg_inst_Result_3_1
    );
  OVtpg_inst_Mcount_Row_cy_3_Q : MUXCY
    port map (
      CI => OVtpg_inst_Mcount_Row_cy(2),
      DI => NlwRenamedSig_OI_vid_field_id,
      S => OVtpg_inst_Mcount_Row_cy_3_rt_319,
      O => OVtpg_inst_Mcount_Row_cy(3)
    );
  OVtpg_inst_Mcount_Row_xor_2_Q : XORCY
    port map (
      CI => OVtpg_inst_Mcount_Row_cy(1),
      LI => OVtpg_inst_Mcount_Row_cy_2_rt_320,
      O => OVtpg_inst_Result_2_1
    );
  OVtpg_inst_Mcount_Row_cy_2_Q : MUXCY
    port map (
      CI => OVtpg_inst_Mcount_Row_cy(1),
      DI => NlwRenamedSig_OI_vid_field_id,
      S => OVtpg_inst_Mcount_Row_cy_2_rt_320,
      O => OVtpg_inst_Mcount_Row_cy(2)
    );
  OVtpg_inst_Mcount_Row_xor_1_Q : XORCY
    port map (
      CI => OVtpg_inst_Mcount_Row_cy(0),
      LI => OVtpg_inst_Mcount_Row_cy_1_rt_321,
      O => OVtpg_inst_Result_1_2
    );
  OVtpg_inst_Mcount_Row_cy_1_Q : MUXCY
    port map (
      CI => OVtpg_inst_Mcount_Row_cy(0),
      DI => NlwRenamedSig_OI_vid_field_id,
      S => OVtpg_inst_Mcount_Row_cy_1_rt_321,
      O => OVtpg_inst_Mcount_Row_cy(1)
    );
  OVtpg_inst_Mcount_Row_xor_0_Q : XORCY
    port map (
      CI => NlwRenamedSig_OI_vid_field_id,
      LI => OVtpg_inst_Mcount_Row_lut(0),
      O => OVtpg_inst_Result_0_2
    );
  OVtpg_inst_Mcount_Row_cy_0_Q : MUXCY
    port map (
      CI => NlwRenamedSig_OI_vid_field_id,
      DI => N1,
      S => OVtpg_inst_Mcount_Row_lut(0),
      O => OVtpg_inst_Mcount_Row_cy(0)
    );
  OVtpg_inst_Mcount_addr_xor_16_Q : XORCY
    port map (
      CI => OVtpg_inst_Mcount_addr_cy(15),
      LI => NlwRenamedSig_OI_OVtpg_inst_addr(16),
      O => OVtpg_inst_Result(16)
    );
  OVtpg_inst_Mcount_addr_xor_15_Q : XORCY
    port map (
      CI => OVtpg_inst_Mcount_addr_cy(14),
      LI => OVtpg_inst_Mcount_addr_cy_15_rt_322,
      O => OVtpg_inst_Result(15)
    );
  OVtpg_inst_Mcount_addr_cy_15_Q : MUXCY
    port map (
      CI => OVtpg_inst_Mcount_addr_cy(14),
      DI => NlwRenamedSig_OI_vid_field_id,
      S => OVtpg_inst_Mcount_addr_cy_15_rt_322,
      O => OVtpg_inst_Mcount_addr_cy(15)
    );
  OVtpg_inst_Mcount_addr_xor_14_Q : XORCY
    port map (
      CI => OVtpg_inst_Mcount_addr_cy(13),
      LI => OVtpg_inst_Mcount_addr_cy_14_rt_323,
      O => OVtpg_inst_Result(14)
    );
  OVtpg_inst_Mcount_addr_cy_14_Q : MUXCY
    port map (
      CI => OVtpg_inst_Mcount_addr_cy(13),
      DI => NlwRenamedSig_OI_vid_field_id,
      S => OVtpg_inst_Mcount_addr_cy_14_rt_323,
      O => OVtpg_inst_Mcount_addr_cy(14)
    );
  OVtpg_inst_Mcount_addr_xor_13_Q : XORCY
    port map (
      CI => OVtpg_inst_Mcount_addr_cy(12),
      LI => OVtpg_inst_Mcount_addr_cy_13_rt_324,
      O => OVtpg_inst_Result(13)
    );
  OVtpg_inst_Mcount_addr_cy_13_Q : MUXCY
    port map (
      CI => OVtpg_inst_Mcount_addr_cy(12),
      DI => NlwRenamedSig_OI_vid_field_id,
      S => OVtpg_inst_Mcount_addr_cy_13_rt_324,
      O => OVtpg_inst_Mcount_addr_cy(13)
    );
  OVtpg_inst_Mcount_addr_xor_12_Q : XORCY
    port map (
      CI => OVtpg_inst_Mcount_addr_cy(11),
      LI => OVtpg_inst_Mcount_addr_cy_12_rt_325,
      O => OVtpg_inst_Result(12)
    );
  OVtpg_inst_Mcount_addr_cy_12_Q : MUXCY
    port map (
      CI => OVtpg_inst_Mcount_addr_cy(11),
      DI => NlwRenamedSig_OI_vid_field_id,
      S => OVtpg_inst_Mcount_addr_cy_12_rt_325,
      O => OVtpg_inst_Mcount_addr_cy(12)
    );
  OVtpg_inst_Mcount_addr_xor_11_Q : XORCY
    port map (
      CI => OVtpg_inst_Mcount_addr_cy(10),
      LI => OVtpg_inst_Mcount_addr_cy_11_rt_326,
      O => OVtpg_inst_Result(11)
    );
  OVtpg_inst_Mcount_addr_cy_11_Q : MUXCY
    port map (
      CI => OVtpg_inst_Mcount_addr_cy(10),
      DI => NlwRenamedSig_OI_vid_field_id,
      S => OVtpg_inst_Mcount_addr_cy_11_rt_326,
      O => OVtpg_inst_Mcount_addr_cy(11)
    );
  OVtpg_inst_Mcount_addr_xor_10_Q : XORCY
    port map (
      CI => OVtpg_inst_Mcount_addr_cy(9),
      LI => OVtpg_inst_Mcount_addr_cy_10_rt_327,
      O => OVtpg_inst_Result(10)
    );
  OVtpg_inst_Mcount_addr_cy_10_Q : MUXCY
    port map (
      CI => OVtpg_inst_Mcount_addr_cy(9),
      DI => NlwRenamedSig_OI_vid_field_id,
      S => OVtpg_inst_Mcount_addr_cy_10_rt_327,
      O => OVtpg_inst_Mcount_addr_cy(10)
    );
  OVtpg_inst_Mcount_addr_xor_9_Q : XORCY
    port map (
      CI => OVtpg_inst_Mcount_addr_cy(8),
      LI => OVtpg_inst_Mcount_addr_cy_9_rt_328,
      O => OVtpg_inst_Result(9)
    );
  OVtpg_inst_Mcount_addr_cy_9_Q : MUXCY
    port map (
      CI => OVtpg_inst_Mcount_addr_cy(8),
      DI => NlwRenamedSig_OI_vid_field_id,
      S => OVtpg_inst_Mcount_addr_cy_9_rt_328,
      O => OVtpg_inst_Mcount_addr_cy(9)
    );
  OVtpg_inst_Mcount_addr_xor_8_Q : XORCY
    port map (
      CI => OVtpg_inst_Mcount_addr_cy(7),
      LI => OVtpg_inst_Mcount_addr_cy_8_rt_329,
      O => OVtpg_inst_Result(8)
    );
  OVtpg_inst_Mcount_addr_cy_8_Q : MUXCY
    port map (
      CI => OVtpg_inst_Mcount_addr_cy(7),
      DI => NlwRenamedSig_OI_vid_field_id,
      S => OVtpg_inst_Mcount_addr_cy_8_rt_329,
      O => OVtpg_inst_Mcount_addr_cy(8)
    );
  OVtpg_inst_Mcount_addr_xor_7_Q : XORCY
    port map (
      CI => OVtpg_inst_Mcount_addr_cy(6),
      LI => OVtpg_inst_Mcount_addr_cy_7_rt_330,
      O => OVtpg_inst_Result(7)
    );
  OVtpg_inst_Mcount_addr_cy_7_Q : MUXCY
    port map (
      CI => OVtpg_inst_Mcount_addr_cy(6),
      DI => NlwRenamedSig_OI_vid_field_id,
      S => OVtpg_inst_Mcount_addr_cy_7_rt_330,
      O => OVtpg_inst_Mcount_addr_cy(7)
    );
  OVtpg_inst_Mcount_addr_xor_6_Q : XORCY
    port map (
      CI => OVtpg_inst_Mcount_addr_cy(5),
      LI => OVtpg_inst_Mcount_addr_cy_6_rt_331,
      O => OVtpg_inst_Result(6)
    );
  OVtpg_inst_Mcount_addr_cy_6_Q : MUXCY
    port map (
      CI => OVtpg_inst_Mcount_addr_cy(5),
      DI => NlwRenamedSig_OI_vid_field_id,
      S => OVtpg_inst_Mcount_addr_cy_6_rt_331,
      O => OVtpg_inst_Mcount_addr_cy(6)
    );
  OVtpg_inst_Mcount_addr_xor_5_Q : XORCY
    port map (
      CI => OVtpg_inst_Mcount_addr_cy(4),
      LI => OVtpg_inst_Mcount_addr_cy_5_rt_332,
      O => OVtpg_inst_Result(5)
    );
  OVtpg_inst_Mcount_addr_cy_5_Q : MUXCY
    port map (
      CI => OVtpg_inst_Mcount_addr_cy(4),
      DI => NlwRenamedSig_OI_vid_field_id,
      S => OVtpg_inst_Mcount_addr_cy_5_rt_332,
      O => OVtpg_inst_Mcount_addr_cy(5)
    );
  OVtpg_inst_Mcount_addr_xor_4_Q : XORCY
    port map (
      CI => OVtpg_inst_Mcount_addr_cy(3),
      LI => OVtpg_inst_Mcount_addr_cy_4_rt_333,
      O => OVtpg_inst_Result(4)
    );
  OVtpg_inst_Mcount_addr_cy_4_Q : MUXCY
    port map (
      CI => OVtpg_inst_Mcount_addr_cy(3),
      DI => NlwRenamedSig_OI_vid_field_id,
      S => OVtpg_inst_Mcount_addr_cy_4_rt_333,
      O => OVtpg_inst_Mcount_addr_cy(4)
    );
  OVtpg_inst_Mcount_addr_xor_3_Q : XORCY
    port map (
      CI => OVtpg_inst_Mcount_addr_cy(2),
      LI => OVtpg_inst_Mcount_addr_cy_3_rt_334,
      O => OVtpg_inst_Result(3)
    );
  OVtpg_inst_Mcount_addr_cy_3_Q : MUXCY
    port map (
      CI => OVtpg_inst_Mcount_addr_cy(2),
      DI => NlwRenamedSig_OI_vid_field_id,
      S => OVtpg_inst_Mcount_addr_cy_3_rt_334,
      O => OVtpg_inst_Mcount_addr_cy(3)
    );
  OVtpg_inst_Mcount_addr_xor_2_Q : XORCY
    port map (
      CI => OVtpg_inst_Mcount_addr_cy(1),
      LI => OVtpg_inst_Mcount_addr_cy_2_rt_335,
      O => OVtpg_inst_Result(2)
    );
  OVtpg_inst_Mcount_addr_cy_2_Q : MUXCY
    port map (
      CI => OVtpg_inst_Mcount_addr_cy(1),
      DI => NlwRenamedSig_OI_vid_field_id,
      S => OVtpg_inst_Mcount_addr_cy_2_rt_335,
      O => OVtpg_inst_Mcount_addr_cy(2)
    );
  OVtpg_inst_Mcount_addr_xor_1_Q : XORCY
    port map (
      CI => OVtpg_inst_Mcount_addr_cy(0),
      LI => OVtpg_inst_Mcount_addr_cy_1_rt_336,
      O => OVtpg_inst_Result_1_1
    );
  OVtpg_inst_Mcount_addr_cy_1_Q : MUXCY
    port map (
      CI => OVtpg_inst_Mcount_addr_cy(0),
      DI => NlwRenamedSig_OI_vid_field_id,
      S => OVtpg_inst_Mcount_addr_cy_1_rt_336,
      O => OVtpg_inst_Mcount_addr_cy(1)
    );
  OVtpg_inst_Mcount_addr_xor_0_Q : XORCY
    port map (
      CI => NlwRenamedSig_OI_vid_field_id,
      LI => OVtpg_inst_Mcount_addr_lut(0),
      O => OVtpg_inst_Result_0_1
    );
  OVtpg_inst_Mcount_addr_cy_0_Q : MUXCY
    port map (
      CI => NlwRenamedSig_OI_vid_field_id,
      DI => N1,
      S => OVtpg_inst_Mcount_addr_lut(0),
      O => OVtpg_inst_Mcount_addr_cy(0)
    );
  OVtpg_inst_Col_10 : FDRE
    port map (
      C => clk_in_100,
      CE => OVtpg_inst_Cen,
      D => OVtpg_inst_Result_10_2,
      R => OVtpg_inst_Mcount_Col_val,
      Q => OVtpg_inst_Col(10)
    );
  OVtpg_inst_Row_10 : FDRE
    port map (
      C => clk_in_100,
      CE => OVtpg_inst_n0315_inv1,
      D => OVtpg_inst_Result_10_1,
      R => OVtpg_inst_Mcount_Row_val,
      Q => OVtpg_inst_Row(10)
    );
  OVtpg_inst_Col_9 : FDRE
    port map (
      C => clk_in_100,
      CE => OVtpg_inst_Cen,
      D => OVtpg_inst_Result_9_2,
      R => OVtpg_inst_Mcount_Col_val,
      Q => OVtpg_inst_Col(9)
    );
  OVtpg_inst_Col_8 : FDRE
    port map (
      C => clk_in_100,
      CE => OVtpg_inst_Cen,
      D => OVtpg_inst_Result_8_2,
      R => OVtpg_inst_Mcount_Col_val,
      Q => OVtpg_inst_Col(8)
    );
  OVtpg_inst_Col_7 : FDRE
    port map (
      C => clk_in_100,
      CE => OVtpg_inst_Cen,
      D => OVtpg_inst_Result_7_2,
      R => OVtpg_inst_Mcount_Col_val,
      Q => OVtpg_inst_Col(7)
    );
  OVtpg_inst_Col_6 : FDRE
    port map (
      C => clk_in_100,
      CE => OVtpg_inst_Cen,
      D => OVtpg_inst_Result_6_2,
      R => OVtpg_inst_Mcount_Col_val,
      Q => OVtpg_inst_Col(6)
    );
  OVtpg_inst_Col_5 : FDRE
    port map (
      C => clk_in_100,
      CE => OVtpg_inst_Cen,
      D => OVtpg_inst_Result_5_2,
      R => OVtpg_inst_Mcount_Col_val,
      Q => OVtpg_inst_Col(5)
    );
  OVtpg_inst_Col_4 : FDRE
    port map (
      C => clk_in_100,
      CE => OVtpg_inst_Cen,
      D => OVtpg_inst_Result_4_2,
      R => OVtpg_inst_Mcount_Col_val,
      Q => OVtpg_inst_Col(4)
    );
  OVtpg_inst_Col_3 : FDRE
    port map (
      C => clk_in_100,
      CE => OVtpg_inst_Cen,
      D => OVtpg_inst_Result_3_2,
      R => OVtpg_inst_Mcount_Col_val,
      Q => OVtpg_inst_Col(3)
    );
  OVtpg_inst_Col_2 : FDRE
    port map (
      C => clk_in_100,
      CE => OVtpg_inst_Cen,
      D => OVtpg_inst_Result_2_2,
      R => OVtpg_inst_Mcount_Col_val,
      Q => OVtpg_inst_Col(2)
    );
  OVtpg_inst_Col_1 : FDRE
    port map (
      C => clk_in_100,
      CE => OVtpg_inst_Cen,
      D => OVtpg_inst_Result_1_3,
      R => OVtpg_inst_Mcount_Col_val,
      Q => OVtpg_inst_Col(1)
    );
  OVtpg_inst_Col_0 : FDRE
    port map (
      C => clk_in_100,
      CE => OVtpg_inst_Cen,
      D => OVtpg_inst_Result_0_3,
      R => OVtpg_inst_Mcount_Col_val,
      Q => OVtpg_inst_Col(0)
    );
  OVtpg_inst_Row_9 : FDRE
    port map (
      C => clk_in_100,
      CE => OVtpg_inst_n0315_inv1,
      D => OVtpg_inst_Result_9_1,
      R => OVtpg_inst_Mcount_Row_val,
      Q => OVtpg_inst_Row(9)
    );
  OVtpg_inst_Row_8 : FDRE
    port map (
      C => clk_in_100,
      CE => OVtpg_inst_n0315_inv1,
      D => OVtpg_inst_Result_8_1,
      R => OVtpg_inst_Mcount_Row_val,
      Q => OVtpg_inst_Row(8)
    );
  OVtpg_inst_Row_7 : FDRE
    port map (
      C => clk_in_100,
      CE => OVtpg_inst_n0315_inv1,
      D => OVtpg_inst_Result_7_1,
      R => OVtpg_inst_Mcount_Row_val,
      Q => OVtpg_inst_Row(7)
    );
  OVtpg_inst_Row_6 : FDRE
    port map (
      C => clk_in_100,
      CE => OVtpg_inst_n0315_inv1,
      D => OVtpg_inst_Result_6_1,
      R => OVtpg_inst_Mcount_Row_val,
      Q => OVtpg_inst_Row(6)
    );
  OVtpg_inst_Row_5 : FDRE
    port map (
      C => clk_in_100,
      CE => OVtpg_inst_n0315_inv1,
      D => OVtpg_inst_Result_5_1,
      R => OVtpg_inst_Mcount_Row_val,
      Q => OVtpg_inst_Row(5)
    );
  OVtpg_inst_Row_4 : FDRE
    port map (
      C => clk_in_100,
      CE => OVtpg_inst_n0315_inv1,
      D => OVtpg_inst_Result_4_1,
      R => OVtpg_inst_Mcount_Row_val,
      Q => OVtpg_inst_Row(4)
    );
  OVtpg_inst_Row_3 : FDRE
    port map (
      C => clk_in_100,
      CE => OVtpg_inst_n0315_inv1,
      D => OVtpg_inst_Result_3_1,
      R => OVtpg_inst_Mcount_Row_val,
      Q => OVtpg_inst_Row(3)
    );
  OVtpg_inst_Row_2 : FDRE
    port map (
      C => clk_in_100,
      CE => OVtpg_inst_n0315_inv1,
      D => OVtpg_inst_Result_2_1,
      R => OVtpg_inst_Mcount_Row_val,
      Q => OVtpg_inst_Row(2)
    );
  OVtpg_inst_Row_1 : FDRE
    port map (
      C => clk_in_100,
      CE => OVtpg_inst_n0315_inv1,
      D => OVtpg_inst_Result_1_2,
      R => OVtpg_inst_Mcount_Row_val,
      Q => OVtpg_inst_Row(1)
    );
  OVtpg_inst_Row_0 : FDRE
    port map (
      C => clk_in_100,
      CE => OVtpg_inst_n0315_inv1,
      D => OVtpg_inst_Result_0_2,
      R => OVtpg_inst_Mcount_Row_val,
      Q => OVtpg_inst_Row(0)
    );
  OVtpg_inst_addr_16 : FDRE
    port map (
      C => clk_in_100,
      CE => OVtpg_inst_n0395_inv,
      D => OVtpg_inst_Result(16),
      R => OVtpg_inst_Mcount_Row_val,
      Q => NlwRenamedSig_OI_OVtpg_inst_addr(16)
    );
  OVtpg_inst_addr_15 : FDRE
    port map (
      C => clk_in_100,
      CE => OVtpg_inst_n0395_inv,
      D => OVtpg_inst_Result(15),
      R => OVtpg_inst_Mcount_Row_val,
      Q => NlwRenamedSig_OI_OVtpg_inst_addr(15)
    );
  OVtpg_inst_addr_14 : FDRE
    port map (
      C => clk_in_100,
      CE => OVtpg_inst_n0395_inv,
      D => OVtpg_inst_Result(14),
      R => OVtpg_inst_Mcount_Row_val,
      Q => NlwRenamedSig_OI_OVtpg_inst_addr(14)
    );
  OVtpg_inst_addr_13 : FDRE
    port map (
      C => clk_in_100,
      CE => OVtpg_inst_n0395_inv,
      D => OVtpg_inst_Result(13),
      R => OVtpg_inst_Mcount_Row_val,
      Q => NlwRenamedSig_OI_OVtpg_inst_addr(13)
    );
  OVtpg_inst_addr_12 : FDRE
    port map (
      C => clk_in_100,
      CE => OVtpg_inst_n0395_inv,
      D => OVtpg_inst_Result(12),
      R => OVtpg_inst_Mcount_Row_val,
      Q => NlwRenamedSig_OI_OVtpg_inst_addr(12)
    );
  OVtpg_inst_addr_11 : FDRE
    port map (
      C => clk_in_100,
      CE => OVtpg_inst_n0395_inv,
      D => OVtpg_inst_Result(11),
      R => OVtpg_inst_Mcount_Row_val,
      Q => NlwRenamedSig_OI_OVtpg_inst_addr(11)
    );
  OVtpg_inst_addr_10 : FDRE
    port map (
      C => clk_in_100,
      CE => OVtpg_inst_n0395_inv,
      D => OVtpg_inst_Result(10),
      R => OVtpg_inst_Mcount_Row_val,
      Q => NlwRenamedSig_OI_OVtpg_inst_addr(10)
    );
  OVtpg_inst_addr_8 : FDRE
    port map (
      C => clk_in_100,
      CE => OVtpg_inst_n0395_inv,
      D => OVtpg_inst_Result(8),
      R => OVtpg_inst_Mcount_Row_val,
      Q => NlwRenamedSig_OI_OVtpg_inst_addr(8)
    );
  OVtpg_inst_addr_7 : FDRE
    port map (
      C => clk_in_100,
      CE => OVtpg_inst_n0395_inv,
      D => OVtpg_inst_Result(7),
      R => OVtpg_inst_Mcount_Row_val,
      Q => NlwRenamedSig_OI_OVtpg_inst_addr(7)
    );
  OVtpg_inst_addr_9 : FDRE
    port map (
      C => clk_in_100,
      CE => OVtpg_inst_n0395_inv,
      D => OVtpg_inst_Result(9),
      R => OVtpg_inst_Mcount_Row_val,
      Q => NlwRenamedSig_OI_OVtpg_inst_addr(9)
    );
  OVtpg_inst_addr_6 : FDRE
    port map (
      C => clk_in_100,
      CE => OVtpg_inst_n0395_inv,
      D => OVtpg_inst_Result(6),
      R => OVtpg_inst_Mcount_Row_val,
      Q => NlwRenamedSig_OI_OVtpg_inst_addr(6)
    );
  OVtpg_inst_addr_5 : FDRE
    port map (
      C => clk_in_100,
      CE => OVtpg_inst_n0395_inv,
      D => OVtpg_inst_Result(5),
      R => OVtpg_inst_Mcount_Row_val,
      Q => NlwRenamedSig_OI_OVtpg_inst_addr(5)
    );
  OVtpg_inst_addr_4 : FDRE
    port map (
      C => clk_in_100,
      CE => OVtpg_inst_n0395_inv,
      D => OVtpg_inst_Result(4),
      R => OVtpg_inst_Mcount_Row_val,
      Q => NlwRenamedSig_OI_OVtpg_inst_addr(4)
    );
  OVtpg_inst_addr_3 : FDRE
    port map (
      C => clk_in_100,
      CE => OVtpg_inst_n0395_inv,
      D => OVtpg_inst_Result(3),
      R => OVtpg_inst_Mcount_Row_val,
      Q => NlwRenamedSig_OI_OVtpg_inst_addr(3)
    );
  OVtpg_inst_addr_2 : FDRE
    port map (
      C => clk_in_100,
      CE => OVtpg_inst_n0395_inv,
      D => OVtpg_inst_Result(2),
      R => OVtpg_inst_Mcount_Row_val,
      Q => NlwRenamedSig_OI_OVtpg_inst_addr(2)
    );
  OVtpg_inst_addr_1 : FDRE
    port map (
      C => clk_in_100,
      CE => OVtpg_inst_n0395_inv,
      D => OVtpg_inst_Result_1_1,
      R => OVtpg_inst_Mcount_Row_val,
      Q => NlwRenamedSig_OI_OVtpg_inst_addr(1)
    );
  OVtpg_inst_addr_0 : FDRE
    port map (
      C => clk_in_100,
      CE => OVtpg_inst_n0395_inv,
      D => OVtpg_inst_Result_0_1,
      R => OVtpg_inst_Mcount_Row_val,
      Q => NlwRenamedSig_OI_OVtpg_inst_addr(0)
    );
  OVtpg_inst_ClkDiv_1 : FDR
    generic map(
      INIT => '0'
    )
    port map (
      C => clk_in_100,
      D => OVtpg_inst_Result(1),
      R => MRST,
      Q => OVtpg_inst_ClkDiv(1)
    );
  OVtpg_inst_ClkDiv_0 : FDR
    generic map(
      INIT => '0'
    )
    port map (
      C => clk_in_100,
      D => OVtpg_inst_PCLK,
      R => MRST,
      Q => OVtpg_inst_ClkDiv(0)
    );
  OVtpg_inst_pmode_2 : FDSE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk_in_100,
      CE => OVtpg_inst_n02371,
      D => OVtpg_inst_Mram_MODE_3_PWR_7_o_wide_mux_9_OUT2,
      S => MRST,
      Q => OVtpg_inst_pmode(2)
    );
  OVtpg_inst_pmode_1 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk_in_100,
      CE => OVtpg_inst_n02371,
      D => OVtpg_inst_Mram_MODE_3_PWR_7_o_wide_mux_9_OUT1,
      R => MRST,
      Q => OVtpg_inst_pmode(1)
    );
  OVtpg_inst_pmode_0 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk_in_100,
      CE => OVtpg_inst_n02371,
      D => OVtpg_inst_Mram_MODE_3_PWR_7_o_wide_mux_9_OUT,
      R => MRST,
      Q => OVtpg_inst_pmode(0)
    );
  OVtpg_inst_HREF : FDE
    port map (
      C => clk_in_100,
      CE => OVtpg_inst_PCLK,
      D => OVtpg_inst_Hrefi_236,
      Q => OVtpg_inst_HREF_61
    );
  OVtpg_inst_VSYNC : FDE
    port map (
      C => clk_in_100,
      CE => OVtpg_inst_PCLK,
      D => OVtpg_inst_Vsynci_237,
      Q => OVtpg_inst_VSYNC_60
    );
  OVtpg_inst_D_7 : FDRE
    port map (
      C => clk_in_100,
      CE => OVtpg_inst_PCLK,
      D => OVtpg_inst_pixel_out_12_pixel_out_23_mux_50_OUT_7_Q,
      R => OVtpg_inst_n0270,
      Q => OVtpg_inst_D(7)
    );
  OVtpg_inst_D_6 : FDRE
    port map (
      C => clk_in_100,
      CE => OVtpg_inst_PCLK,
      D => OVtpg_inst_pixel_out_12_pixel_out_23_mux_50_OUT_6_Q,
      R => OVtpg_inst_n0270,
      Q => OVtpg_inst_D(6)
    );
  OVtpg_inst_D_5 : FDRE
    port map (
      C => clk_in_100,
      CE => OVtpg_inst_PCLK,
      D => OVtpg_inst_pixel_out_12_pixel_out_23_mux_50_OUT_5_Q,
      R => OVtpg_inst_n0270,
      Q => OVtpg_inst_D(5)
    );
  OVtpg_inst_D_4 : FDRE
    port map (
      C => clk_in_100,
      CE => OVtpg_inst_PCLK,
      D => OVtpg_inst_pixel_out_12_pixel_out_23_mux_50_OUT_4_Q,
      R => OVtpg_inst_n0270,
      Q => OVtpg_inst_D(4)
    );
  OVtpg_inst_D_3 : FDRE
    port map (
      C => clk_in_100,
      CE => OVtpg_inst_PCLK,
      D => OVtpg_inst_pixel_out_12_pixel_out_23_mux_50_OUT_3_Q,
      R => OVtpg_inst_n0270,
      Q => OVtpg_inst_D(3)
    );
  OVtpg_inst_D_2 : FDRE
    port map (
      C => clk_in_100,
      CE => OVtpg_inst_PCLK,
      D => OVtpg_inst_pixel_out_12_pixel_out_23_mux_50_OUT_2_Q,
      R => OVtpg_inst_n0270,
      Q => OVtpg_inst_D(2)
    );
  OVtpg_inst_D_1 : FDRE
    port map (
      C => clk_in_100,
      CE => OVtpg_inst_PCLK,
      D => OVtpg_inst_pixel_out_12_pixel_out_23_mux_50_OUT_1_Q,
      R => OVtpg_inst_n0270,
      Q => OVtpg_inst_D(1)
    );
  OVtpg_inst_D_0 : FDRE
    port map (
      C => clk_in_100,
      CE => OVtpg_inst_PCLK,
      D => OVtpg_inst_pixel_out_12_pixel_out_23_mux_50_OUT_0_Q,
      R => OVtpg_inst_n0270,
      Q => OVtpg_inst_D(0)
    );
  SIF_inst_RGB_data_23 : FDRE
    port map (
      C => clk_in_50,
      CE => SIF_inst_oddpix1,
      D => SIF_inst_FirstByte(7),
      R => SIF_inst_Reset_OR_DriverANDClockEnable,
      Q => NlwRenamedSignal_SIF_inst_RGB_data_23_Q
    );
  SIF_inst_RGB_data_22 : FDRE
    port map (
      C => clk_in_50,
      CE => SIF_inst_oddpix1,
      D => SIF_inst_FirstByte(6),
      R => SIF_inst_Reset_OR_DriverANDClockEnable,
      Q => NlwRenamedSignal_SIF_inst_RGB_data_22_Q
    );
  SIF_inst_RGB_data_21 : FDRE
    port map (
      C => clk_in_50,
      CE => SIF_inst_oddpix1,
      D => SIF_inst_FirstByte(5),
      R => SIF_inst_Reset_OR_DriverANDClockEnable,
      Q => NlwRenamedSignal_SIF_inst_RGB_data_21_Q
    );
  SIF_inst_RGB_data_20 : FDRE
    port map (
      C => clk_in_50,
      CE => SIF_inst_oddpix1,
      D => SIF_inst_FirstByte(4),
      R => SIF_inst_Reset_OR_DriverANDClockEnable,
      Q => NlwRenamedSignal_SIF_inst_RGB_data_20_Q
    );
  SIF_inst_RGB_data_16 : FDRE
    port map (
      C => clk_in_50,
      CE => SIF_inst_oddpix1,
      D => SIF_inst_FirstByte(3),
      R => SIF_inst_Reset_OR_DriverANDClockEnable,
      Q => NlwRenamedSignal_SIF_inst_RGB_data_16_Q
    );
  SIF_inst_RGB_data_15 : FDRE
    port map (
      C => clk_in_50,
      CE => SIF_inst_oddpix1,
      D => SIF_inst_FirstByte(2),
      R => SIF_inst_Reset_OR_DriverANDClockEnable,
      Q => NlwRenamedSignal_SIF_inst_RGB_data_15_Q
    );
  SIF_inst_RGB_data_14 : FDRE
    port map (
      C => clk_in_50,
      CE => SIF_inst_oddpix1,
      D => SIF_inst_FirstByte(1),
      R => SIF_inst_Reset_OR_DriverANDClockEnable,
      Q => NlwRenamedSignal_SIF_inst_RGB_data_14_Q
    );
  SIF_inst_RGB_data_13 : FDRE
    port map (
      C => clk_in_50,
      CE => SIF_inst_oddpix1,
      D => SIF_inst_FirstByte(0),
      R => SIF_inst_Reset_OR_DriverANDClockEnable,
      Q => NlwRenamedSignal_SIF_inst_RGB_data_13_Q
    );
  SIF_inst_RGB_data_12 : FDRE
    port map (
      C => clk_in_50,
      CE => SIF_inst_oddpix1,
      D => OVtpg_inst_D(7),
      R => SIF_inst_Reset_OR_DriverANDClockEnable,
      Q => NlwRenamedSignal_SIF_inst_RGB_data_12_Q
    );
  SIF_inst_RGB_data_11 : FDRE
    port map (
      C => clk_in_50,
      CE => SIF_inst_oddpix1,
      D => OVtpg_inst_D(6),
      R => SIF_inst_Reset_OR_DriverANDClockEnable,
      Q => NlwRenamedSignal_SIF_inst_RGB_data_11_Q
    );
  SIF_inst_RGB_data_8 : FDRE
    port map (
      C => clk_in_50,
      CE => SIF_inst_oddpix1,
      D => OVtpg_inst_D(5),
      R => SIF_inst_Reset_OR_DriverANDClockEnable,
      Q => NlwRenamedSignal_SIF_inst_RGB_data_8_Q
    );
  SIF_inst_RGB_data_7 : FDRE
    port map (
      C => clk_in_50,
      CE => SIF_inst_oddpix1,
      D => OVtpg_inst_D(4),
      R => SIF_inst_Reset_OR_DriverANDClockEnable,
      Q => NlwRenamedSignal_SIF_inst_RGB_data_7_Q
    );
  SIF_inst_RGB_data_6 : FDRE
    port map (
      C => clk_in_50,
      CE => SIF_inst_oddpix1,
      D => OVtpg_inst_D(3),
      R => SIF_inst_Reset_OR_DriverANDClockEnable,
      Q => NlwRenamedSignal_SIF_inst_RGB_data_6_Q
    );
  SIF_inst_RGB_data_5 : FDRE
    port map (
      C => clk_in_50,
      CE => SIF_inst_oddpix1,
      D => OVtpg_inst_D(2),
      R => SIF_inst_Reset_OR_DriverANDClockEnable,
      Q => NlwRenamedSignal_SIF_inst_RGB_data_5_Q
    );
  SIF_inst_RGB_data_4 : FDRE
    port map (
      C => clk_in_50,
      CE => SIF_inst_oddpix1,
      D => OVtpg_inst_D(1),
      R => SIF_inst_Reset_OR_DriverANDClockEnable,
      Q => NlwRenamedSignal_SIF_inst_RGB_data_4_Q
    );
  SIF_inst_RGB_data_0 : FDRE
    port map (
      C => clk_in_50,
      CE => SIF_inst_oddpix1,
      D => OVtpg_inst_D(0),
      R => SIF_inst_Reset_OR_DriverANDClockEnable,
      Q => NlwRenamedSignal_SIF_inst_RGB_data_0_Q
    );
  SIF_inst_Vsync : FDSE
    port map (
      C => clk_in_50,
      CE => SIF_inst_oddpix1,
      D => SIF_inst_VS_in_INV_360_o,
      S => MRST,
      Q => NlwRenamedSig_OI_SIF_inst_Vsync
    );
  SIF_inst_Hsync : FDSE
    port map (
      C => clk_in_50,
      CE => SIF_inst_oddpix1,
      D => OVtpg_inst_Hsynci_234,
      S => MRST,
      Q => NlwRenamedSig_OI_SIF_inst_Hsync
    );
  SIF_inst_oddpix : FDR
    port map (
      C => clk_in_50,
      D => SIF_inst_oddpix_INV_358_o,
      R => SIF_inst_Reset_OR_DriverANDClockEnable,
      Q => SIF_inst_oddpix_252
    );
  SIF_inst_FirstByte_7 : FDE
    port map (
      C => clk_in_50,
      CE => SIF_inst_n0060_inv,
      D => OVtpg_inst_D(7),
      Q => SIF_inst_FirstByte(7)
    );
  SIF_inst_FirstByte_6 : FDE
    port map (
      C => clk_in_50,
      CE => SIF_inst_n0060_inv,
      D => OVtpg_inst_D(6),
      Q => SIF_inst_FirstByte(6)
    );
  SIF_inst_FirstByte_5 : FDE
    port map (
      C => clk_in_50,
      CE => SIF_inst_n0060_inv,
      D => OVtpg_inst_D(5),
      Q => SIF_inst_FirstByte(5)
    );
  SIF_inst_FirstByte_4 : FDE
    port map (
      C => clk_in_50,
      CE => SIF_inst_n0060_inv,
      D => OVtpg_inst_D(4),
      Q => SIF_inst_FirstByte(4)
    );
  SIF_inst_FirstByte_3 : FDE
    port map (
      C => clk_in_50,
      CE => SIF_inst_n0060_inv,
      D => OVtpg_inst_D(3),
      Q => SIF_inst_FirstByte(3)
    );
  SIF_inst_FirstByte_2 : FDE
    port map (
      C => clk_in_50,
      CE => SIF_inst_n0060_inv,
      D => OVtpg_inst_D(2),
      Q => SIF_inst_FirstByte(2)
    );
  SIF_inst_FirstByte_1 : FDE
    port map (
      C => clk_in_50,
      CE => SIF_inst_n0060_inv,
      D => OVtpg_inst_D(1),
      Q => SIF_inst_FirstByte(1)
    );
  SIF_inst_FirstByte_0 : FDE
    port map (
      C => clk_in_50,
      CE => SIF_inst_n0060_inv,
      D => OVtpg_inst_D(0),
      Q => SIF_inst_FirstByte(0)
    );
  OVtpg_inst_n023711 : LUT6
    generic map(
      INIT => X"0000000000200000"
    )
    port map (
      I0 => OVtpg_inst_n0315_inv1,
      I1 => OVtpg_inst_Row(1),
      I2 => OVtpg_inst_Row_10_GND_7_o_equal_8_o_10_1,
      I3 => OVtpg_inst_Row(2),
      I4 => OVtpg_inst_Row(5),
      I5 => OVtpg_inst_Row(4),
      O => OVtpg_inst_n02371
    );
  OVtpg_inst_Mmux_pixel_out_12_pixel_out_23_mux_50_OUT31121 : LUT3
    generic map(
      INIT => X"57"
    )
    port map (
      I0 => OVtpg_inst_pmode(0),
      I1 => OVtpg_inst_n0134(3),
      I2 => OVtpg_inst_n0134(2),
      O => OVtpg_inst_Mmux_pixel_out_12_pixel_out_23_mux_50_OUT3112
    );
  OVtpg_inst_Mmux_pixel_out_12_pixel_out_23_mux_50_OUT31421 : LUT4
    generic map(
      INIT => X"EAAA"
    )
    port map (
      I0 => OVtpg_inst_n0134(3),
      I1 => OVtpg_inst_n0134(2),
      I2 => OVtpg_inst_n0134(1),
      I3 => OVtpg_inst_n0134(0),
      O => OVtpg_inst_Mmux_pixel_out_12_pixel_out_23_mux_50_OUT3142
    );
  OVtpg_inst_Mram_MODE_3_PWR_7_o_wide_mux_9_OUT21 : LUT4
    generic map(
      INIT => X"FFE8"
    )
    port map (
      I0 => mode_sel(1),
      I1 => mode_sel(3),
      I2 => mode_sel(0),
      I3 => mode_sel(2),
      O => OVtpg_inst_Mram_MODE_3_PWR_7_o_wide_mux_9_OUT2
    );
  OVtpg_inst_Mram_MODE_3_PWR_7_o_wide_mux_9_OUT111 : LUT4
    generic map(
      INIT => X"0110"
    )
    port map (
      I0 => mode_sel(0),
      I1 => mode_sel(2),
      I2 => mode_sel(1),
      I3 => mode_sel(3),
      O => OVtpg_inst_Mram_MODE_3_PWR_7_o_wide_mux_9_OUT1
    );
  OVtpg_inst_Mram_MODE_3_PWR_7_o_wide_mux_9_OUT11 : LUT4
    generic map(
      INIT => X"0110"
    )
    port map (
      I0 => mode_sel(1),
      I1 => mode_sel(2),
      I2 => mode_sel(0),
      I3 => mode_sel(3),
      O => OVtpg_inst_Mram_MODE_3_PWR_7_o_wide_mux_9_OUT
    );
  OVtpg_inst_Mcount_Row_val1 : LUT6
    generic map(
      INIT => X"555D555555555555"
    )
    port map (
      I0 => locked_in,
      I1 => OVtpg_inst_Row(2),
      I2 => OVtpg_inst_Row(1),
      I3 => OVtpg_inst_Row(0),
      I4 => OVtpg_inst_Row_10_GND_7_o_equal_5_o_10_1_96,
      I5 => OVtpg_inst_n0315_inv1,
      O => OVtpg_inst_Mcount_Row_val
    );
  OVtpg_inst_Col_10_GND_7_o_equal_4_o_10_2 : LUT6
    generic map(
      INIT => X"0002000000000000"
    )
    port map (
      I0 => OVtpg_inst_Col(4),
      I1 => OVtpg_inst_Col(5),
      I2 => OVtpg_inst_Col(6),
      I3 => OVtpg_inst_Col(7),
      I4 => OVtpg_inst_Col(8),
      I5 => OVtpg_inst_Col_10_GND_7_o_equal_4_o_10_1,
      O => OVtpg_inst_Col_10_GND_7_o_equal_4_o
    );
  OVtpg_inst_Col_10_GND_7_o_equal_4_o_10_11 : LUT6
    generic map(
      INIT => X"0000800000000000"
    )
    port map (
      I0 => OVtpg_inst_Col(0),
      I1 => OVtpg_inst_Col(1),
      I2 => OVtpg_inst_Col(2),
      I3 => OVtpg_inst_Col(3),
      I4 => OVtpg_inst_Col(10),
      I5 => OVtpg_inst_Col(9),
      O => OVtpg_inst_Col_10_GND_7_o_equal_4_o_10_1
    );
  OVtpg_inst_n0315_inv11 : LUT3
    generic map(
      INIT => X"80"
    )
    port map (
      I0 => OVtpg_inst_ClkDiv(1),
      I1 => OVtpg_inst_ClkDiv(0),
      I2 => OVtpg_inst_Col_10_GND_7_o_equal_4_o,
      O => OVtpg_inst_n0315_inv1
    );
  OVtpg_inst_Mcount_ClkDiv_xor_1_11 : LUT2
    generic map(
      INIT => X"6"
    )
    port map (
      I0 => OVtpg_inst_ClkDiv(1),
      I1 => OVtpg_inst_ClkDiv(0),
      O => OVtpg_inst_Result(1)
    );
  OVtpg_inst_n02701 : LUT2
    generic map(
      INIT => X"1"
    )
    port map (
      I0 => OVtpg_inst_ClkDiv(0),
      I1 => OVtpg_inst_Hrefi_236,
      O => OVtpg_inst_n0270
    );
  OVtpg_inst_Cen_1_1 : LUT2
    generic map(
      INIT => X"8"
    )
    port map (
      I0 => OVtpg_inst_ClkDiv(1),
      I1 => OVtpg_inst_ClkDiv(0),
      O => OVtpg_inst_Cen
    );
  OVtpg_inst_Row_10_PWR_7_o_div_45_Madd_a_10_GND_9_o_add_17_OUT_10_0_cy_9_11 : LUT6
    generic map(
      INIT => X"787878707870F0F0"
    )
    port map (
      I0 => OVtpg_inst_Row(7),
      I1 => OVtpg_inst_Row(8),
      I2 => OVtpg_inst_Row(9),
      I3 => OVtpg_inst_Row(5),
      I4 => OVtpg_inst_Row(6),
      I5 => OVtpg_inst_Row(10),
      O => OVtpg_inst_n0134(3)
    );
  OVtpg_inst_Col_10_PWR_7_o_div_44_o_0_11 : LUT6
    generic map(
      INIT => X"FFFF380EFFFF83E0"
    )
    port map (
      I0 => OVtpg_inst_Col(4),
      I1 => OVtpg_inst_Col(5),
      I2 => OVtpg_inst_Col(6),
      I3 => OVtpg_inst_Col_10_PWR_7_o_div_44_Madd_a_10_GND_8_o_add_21_OUT_10_0_lut_7_Q,
      I4 => OVtpg_inst_Col_10_PWR_7_o_div_44_o_0_13,
      I5 => OVtpg_inst_n0133(2),
      O => OVtpg_inst_n0133(0)
    );
  OVtpg_inst_Col_10_PWR_7_o_div_44_o_0_131 : LUT5
    generic map(
      INIT => X"10088160"
    )
    port map (
      I0 => OVtpg_inst_Col(6),
      I1 => OVtpg_inst_Col(10),
      I2 => OVtpg_inst_Col(9),
      I3 => OVtpg_inst_Col(8),
      I4 => OVtpg_inst_Col(7),
      O => OVtpg_inst_Col_10_PWR_7_o_div_44_o_0_13
    );
  OVtpg_inst_Col_10_PWR_7_o_div_44_o_2_1 : LUT5
    generic map(
      INIT => X"0BC2F0BC"
    )
    port map (
      I0 => OVtpg_inst_Col(6),
      I1 => OVtpg_inst_Col(9),
      I2 => OVtpg_inst_Col(10),
      I3 => OVtpg_inst_Col(7),
      I4 => OVtpg_inst_Col(8),
      O => OVtpg_inst_n0133(2)
    );
  OVtpg_inst_Col_10_PWR_7_o_div_44_Mmux_n045991 : LUT5
    generic map(
      INIT => X"0E877018"
    )
    port map (
      I0 => OVtpg_inst_Col(6),
      I1 => OVtpg_inst_Col(10),
      I2 => OVtpg_inst_Col(9),
      I3 => OVtpg_inst_Col(8),
      I4 => OVtpg_inst_Col(7),
      O => OVtpg_inst_Col_10_PWR_7_o_div_44_Madd_a_10_GND_8_o_add_21_OUT_10_0_lut_7_Q
    );
  OVtpg_inst_Col_10_PWR_7_o_div_44_o_3_1 : LUT4
    generic map(
      INIT => X"91A8"
    )
    port map (
      I0 => OVtpg_inst_Col(9),
      I1 => OVtpg_inst_Col(8),
      I2 => OVtpg_inst_Col(7),
      I3 => OVtpg_inst_Col(10),
      O => OVtpg_inst_n0133(3)
    );
  SIF_inst_Reset_OR_DriverANDClockEnable491 : LUT2
    generic map(
      INIT => X"7"
    )
    port map (
      I0 => locked_in,
      I1 => OVtpg_inst_HREF_61,
      O => SIF_inst_Reset_OR_DriverANDClockEnable
    );
  SIF_inst_n0060_inv1 : LUT3
    generic map(
      INIT => X"08"
    )
    port map (
      I0 => locked_in,
      I1 => OVtpg_inst_HREF_61,
      I2 => SIF_inst_oddpix_252,
      O => SIF_inst_n0060_inv
    );
  SIF_inst_oddpix11 : LUT2
    generic map(
      INIT => X"B"
    )
    port map (
      I0 => SIF_inst_oddpix_252,
      I1 => OVtpg_inst_HREF_61,
      O => SIF_inst_oddpix1
    );
  OVtpg_inst_Mmux_pixel_out_12_pixel_out_23_mux_50_OUT3173 : LUT6
    generic map(
      INIT => X"5555555554445000"
    )
    port map (
      I0 => OVtpg_inst_pmode(1),
      I1 => OVtpg_inst_Mmux_pixel_out_12_pixel_out_23_mux_50_OUT3172_262,
      I2 => OVtpg_inst_Mmux_pixel_out_12_pixel_out_23_mux_50_OUT3171_261,
      I3 => OVtpg_inst_Mmux_pixel_out_12_pixel_out_23_mux_50_OUT3111,
      I4 => OVtpg_inst_Mmux_pixel_out_12_pixel_out_23_mux_50_OUT3112,
      I5 => OVtpg_inst_Mmux_pixel_out_12_pixel_out_23_mux_50_OUT3113,
      O => OVtpg_inst_Mmux_pixel_out_12_pixel_out_23_mux_50_OUT3173_263
    );
  OVtpg_inst_Mmux_pixel_out_12_pixel_out_23_mux_50_OUT3174 : LUT2
    generic map(
      INIT => X"2"
    )
    port map (
      I0 => OVtpg_inst_pmode(1),
      I1 => OVtpg_inst_pmode(0),
      O => OVtpg_inst_Mmux_pixel_out_12_pixel_out_23_mux_50_OUT3164
    );
  OVtpg_inst_Mmux_pixel_out_12_pixel_out_23_mux_50_OUT3179 : LUT6
    generic map(
      INIT => X"FFFF8A0AFFFF8800"
    )
    port map (
      I0 => OVtpg_inst_Mmux_pixel_out_12_pixel_out_23_mux_50_OUT3164,
      I1 => OVtpg_inst_Mmux_pixel_out_12_pixel_out_23_mux_50_OUT3178_265,
      I2 => OVtpg_inst_n0134(3),
      I3 => OVtpg_inst_Mmux_pixel_out_12_pixel_out_23_mux_50_OUT3142,
      I4 => OVtpg_inst_Mmux_pixel_out_12_pixel_out_23_mux_50_OUT3173_263,
      I5 => OVtpg_inst_Mmux_pixel_out_12_pixel_out_23_mux_50_OUT3177_264,
      O => OVtpg_inst_Mmux_pixel_out_12_pixel_out_23_mux_50_OUT317
    );
  OVtpg_inst_Mmux_pixel_out_12_pixel_out_23_mux_50_OUT41121 : LUT2
    generic map(
      INIT => X"8"
    )
    port map (
      I0 => OVtpg_inst_pmode(0),
      I1 => OVtpg_inst_n0133(1),
      O => OVtpg_inst_Mmux_pixel_out_12_pixel_out_23_mux_50_OUT41121_266
    );
  OVtpg_inst_Mmux_pixel_out_12_pixel_out_23_mux_50_OUT41123 : LUT6
    generic map(
      INIT => X"5555555554445000"
    )
    port map (
      I0 => OVtpg_inst_pmode(1),
      I1 => OVtpg_inst_Mmux_pixel_out_12_pixel_out_23_mux_50_OUT41122_267,
      I2 => OVtpg_inst_Mmux_pixel_out_12_pixel_out_23_mux_50_OUT41121_266,
      I3 => OVtpg_inst_Mmux_pixel_out_12_pixel_out_23_mux_50_OUT3111,
      I4 => OVtpg_inst_Mmux_pixel_out_12_pixel_out_23_mux_50_OUT3112,
      I5 => OVtpg_inst_Mmux_pixel_out_12_pixel_out_23_mux_50_OUT3113,
      O => OVtpg_inst_Mmux_pixel_out_12_pixel_out_23_mux_50_OUT41123_268
    );
  OVtpg_inst_Mmux_pixel_out_12_pixel_out_23_mux_50_OUT41129 : LUT5
    generic map(
      INIT => X"F2F2F2F0"
    )
    port map (
      I0 => OVtpg_inst_pmode(1),
      I1 => OVtpg_inst_pmode(0),
      I2 => OVtpg_inst_Mmux_pixel_out_12_pixel_out_23_mux_50_OUT41123_268,
      I3 => OVtpg_inst_Mmux_pixel_out_12_pixel_out_23_mux_50_OUT41128_271,
      I4 => OVtpg_inst_Mmux_pixel_out_12_pixel_out_23_mux_50_OUT41126_270,
      O => OVtpg_inst_Mmux_pixel_out_12_pixel_out_23_mux_50_OUT4112
    );
  OVtpg_inst_n0358_inv_SW0 : LUT4
    generic map(
      INIT => X"BFFF"
    )
    port map (
      I0 => OVtpg_inst_Col(4),
      I1 => OVtpg_inst_Col(5),
      I2 => OVtpg_inst_ClkDiv(1),
      I3 => OVtpg_inst_ClkDiv(0),
      O => N4
    );
  OVtpg_inst_n0358_inv : LUT6
    generic map(
      INIT => X"0000000000200000"
    )
    port map (
      I0 => OVtpg_inst_Col_10_GND_7_o_equal_4_o_10_1,
      I1 => OVtpg_inst_Col_10_GND_7_o_equal_4_o,
      I2 => OVtpg_inst_Col(7),
      I3 => OVtpg_inst_Col(8),
      I4 => OVtpg_inst_Col(6),
      I5 => N4,
      O => OVtpg_inst_n0358_inv_184
    );
  OVtpg_inst_n0262_SW0 : LUT5
    generic map(
      INIT => X"FFFFBFFF"
    )
    port map (
      I0 => OVtpg_inst_Col(4),
      I1 => OVtpg_inst_ClkDiv(1),
      I2 => OVtpg_inst_ClkDiv(0),
      I3 => locked_in,
      I4 => OVtpg_inst_Col(5),
      O => N6
    );
  OVtpg_inst_n0244_SW0 : LUT5
    generic map(
      INIT => X"80000000"
    )
    port map (
      I0 => OVtpg_inst_Col(5),
      I1 => OVtpg_inst_Col(4),
      I2 => OVtpg_inst_ClkDiv(1),
      I3 => OVtpg_inst_ClkDiv(0),
      I4 => locked_in,
      O => N8
    );
  OVtpg_inst_n0244 : LUT6
    generic map(
      INIT => X"0000000000200000"
    )
    port map (
      I0 => OVtpg_inst_Col_10_GND_7_o_equal_4_o_10_1,
      I1 => OVtpg_inst_Col_10_GND_7_o_equal_4_o,
      I2 => N8,
      I3 => OVtpg_inst_Col(7),
      I4 => OVtpg_inst_Col(6),
      I5 => OVtpg_inst_Col(8),
      O => OVtpg_inst_n0244_198
    );
  OVtpg_inst_n0395_inv4 : LUT5
    generic map(
      INIT => X"08000000"
    )
    port map (
      I0 => OVtpg_inst_n0395_inv3_275,
      I1 => OVtpg_inst_Inside,
      I2 => OVtpg_inst_Col_10_GND_7_o_equal_4_o,
      I3 => OVtpg_inst_ClkDiv(0),
      I4 => OVtpg_inst_ClkDiv(1),
      O => OVtpg_inst_n0395_inv
    );
  OVtpg_inst_Mmux_pixel_out_12_pixel_out_23_mux_50_OUT71 : LUT5
    generic map(
      INIT => X"CCF000AA"
    )
    port map (
      I0 => test_data(10),
      I1 => rom_dat(6),
      I2 => rom_dat(14),
      I3 => OVtpg_inst_ClkDiv(1),
      I4 => OVtpg_inst_Inside,
      O => OVtpg_inst_Mmux_pixel_out_12_pixel_out_23_mux_50_OUT7
    );
  OVtpg_inst_Mmux_pixel_out_12_pixel_out_23_mux_50_OUT72 : LUT4
    generic map(
      INIT => X"EAAA"
    )
    port map (
      I0 => OVtpg_inst_pmode(2),
      I1 => OVtpg_inst_pmode(1),
      I2 => OVtpg_inst_pmode(0),
      I3 => OVtpg_inst_Mmux_pixel_out_12_pixel_out_23_mux_50_OUT7,
      O => OVtpg_inst_Mmux_pixel_out_12_pixel_out_23_mux_50_OUT71_277
    );
  OVtpg_inst_Mmux_pixel_out_12_pixel_out_23_mux_50_OUT61 : LUT5
    generic map(
      INIT => X"CCF000AA"
    )
    port map (
      I0 => test_data(9),
      I1 => rom_dat(5),
      I2 => rom_dat(13),
      I3 => OVtpg_inst_ClkDiv(1),
      I4 => OVtpg_inst_Inside,
      O => OVtpg_inst_Mmux_pixel_out_12_pixel_out_23_mux_50_OUT6
    );
  OVtpg_inst_Mmux_pixel_out_12_pixel_out_23_mux_50_OUT62 : LUT4
    generic map(
      INIT => X"EAAA"
    )
    port map (
      I0 => OVtpg_inst_pmode(2),
      I1 => OVtpg_inst_pmode(1),
      I2 => OVtpg_inst_pmode(0),
      I3 => OVtpg_inst_Mmux_pixel_out_12_pixel_out_23_mux_50_OUT6,
      O => OVtpg_inst_Mmux_pixel_out_12_pixel_out_23_mux_50_OUT61_279
    );
  OVtpg_inst_Mmux_pixel_out_12_pixel_out_23_mux_50_OUT81 : LUT6
    generic map(
      INIT => X"F0F000CC000000AA"
    )
    port map (
      I0 => test_data(11),
      I1 => rom_dat(15),
      I2 => rom_dat(7),
      I3 => OVtpg_inst_pmode(2),
      I4 => OVtpg_inst_ClkDiv(1),
      I5 => OVtpg_inst_Inside,
      O => OVtpg_inst_Mmux_pixel_out_12_pixel_out_23_mux_50_OUT8
    );
  OVtpg_inst_Mmux_pixel_out_12_pixel_out_23_mux_50_OUT2_SW0 : LUT6
    generic map(
      INIT => X"F0F000CC000000AA"
    )
    port map (
      I0 => test_data(6),
      I1 => rom_dat(9),
      I2 => rom_dat(1),
      I3 => OVtpg_inst_pmode(2),
      I4 => OVtpg_inst_ClkDiv(1),
      I5 => OVtpg_inst_Inside,
      O => N10
    );
  OVtpg_inst_Mmux_pixel_out_12_pixel_out_23_mux_50_OUT5_SW0 : LUT6
    generic map(
      INIT => X"FF335555FF0FFFFF"
    )
    port map (
      I0 => rom_dat(12),
      I1 => rom_dat(4),
      I2 => test_data(3),
      I3 => OVtpg_inst_pmode(2),
      I4 => OVtpg_inst_ClkDiv(1),
      I5 => OVtpg_inst_Inside,
      O => N12
    );
  OVtpg_inst_Mmux_pixel_out_12_pixel_out_23_mux_50_OUT4_SW0 : LUT6
    generic map(
      INIT => X"FF335555FF0FFFFF"
    )
    port map (
      I0 => rom_dat(11),
      I1 => rom_dat(3),
      I2 => test_data(2),
      I3 => OVtpg_inst_pmode(2),
      I4 => OVtpg_inst_ClkDiv(1),
      I5 => OVtpg_inst_Inside,
      O => N14
    );
  OVtpg_inst_Mmux_pixel_out_12_pixel_out_23_mux_50_OUT1_SW0 : LUT6
    generic map(
      INIT => X"F0F000CC000000AA"
    )
    port map (
      I0 => test_data(5),
      I1 => rom_dat(8),
      I2 => rom_dat(0),
      I3 => OVtpg_inst_pmode(2),
      I4 => OVtpg_inst_ClkDiv(1),
      I5 => OVtpg_inst_Inside,
      O => N16
    );
  OVtpg_inst_Mmux_pixel_out_12_pixel_out_23_mux_50_OUT31 : LUT6
    generic map(
      INIT => X"F0F0CCCCFF00AAAA"
    )
    port map (
      I0 => test_data(7),
      I1 => rom_dat(10),
      I2 => rom_dat(2),
      I3 => test_data(1),
      I4 => OVtpg_inst_ClkDiv(1),
      I5 => OVtpg_inst_Inside,
      O => OVtpg_inst_Mmux_pixel_out_12_pixel_out_23_mux_50_OUT3
    );
  OVtpg_inst_Mmux_pixel_out_12_pixel_out_23_mux_50_OUT32 : LUT3
    generic map(
      INIT => X"80"
    )
    port map (
      I0 => OVtpg_inst_pmode(1),
      I1 => OVtpg_inst_pmode(0),
      I2 => OVtpg_inst_Mmux_pixel_out_12_pixel_out_23_mux_50_OUT3,
      O => OVtpg_inst_Mmux_pixel_out_12_pixel_out_23_mux_50_OUT31_286
    );
  OVtpg_inst_Mmux_pixel_out_12_pixel_out_23_mux_50_OUT33 : LUT5
    generic map(
      INIT => X"55545150"
    )
    port map (
      I0 => OVtpg_inst_pmode(2),
      I1 => OVtpg_inst_ClkDiv(1),
      I2 => OVtpg_inst_Mmux_pixel_out_12_pixel_out_23_mux_50_OUT31_286,
      I3 => OVtpg_inst_Mmux_pixel_out_12_pixel_out_23_mux_50_OUT317,
      I4 => OVtpg_inst_Mmux_pixel_out_12_pixel_out_23_mux_50_OUT316,
      O => OVtpg_inst_pixel_out_12_pixel_out_23_mux_50_OUT_2_Q
    );
  OVtpg_inst_Inside1 : LUT6
    generic map(
      INIT => X"0F380F700FF00FF0"
    )
    port map (
      I0 => OVtpg_inst_Row(3),
      I1 => OVtpg_inst_Row(6),
      I2 => OVtpg_inst_Row(8),
      I3 => OVtpg_inst_Row(7),
      I4 => OVtpg_inst_Row(4),
      I5 => OVtpg_inst_Row(5),
      O => OVtpg_inst_Inside1_287
    );
  OVtpg_inst_Inside2 : LUT6
    generic map(
      INIT => X"0111101011111000"
    )
    port map (
      I0 => OVtpg_inst_Row(9),
      I1 => OVtpg_inst_Row(10),
      I2 => OVtpg_inst_Col(7),
      I3 => OVtpg_inst_Col(5),
      I4 => OVtpg_inst_Col(8),
      I5 => OVtpg_inst_Col(6),
      O => OVtpg_inst_Inside2_288
    );
  OVtpg_inst_Inside3 : LUT4
    generic map(
      INIT => X"1000"
    )
    port map (
      I0 => OVtpg_inst_Col(9),
      I1 => OVtpg_inst_Col(10),
      I2 => OVtpg_inst_Inside1_287,
      I3 => OVtpg_inst_Inside2_288,
      O => OVtpg_inst_Inside
    );
  OVtpg_inst_n0315_inv2_SW0 : LUT2
    generic map(
      INIT => X"B"
    )
    port map (
      I0 => OVtpg_inst_Row(0),
      I1 => OVtpg_inst_Row(3),
      O => N18
    );
  OVtpg_inst_n0315_inv2 : LUT6
    generic map(
      INIT => X"0000000000200000"
    )
    port map (
      I0 => OVtpg_inst_Row(7),
      I1 => OVtpg_inst_Row(10),
      I2 => OVtpg_inst_Row(8),
      I3 => OVtpg_inst_Row(9),
      I4 => OVtpg_inst_Row(6),
      I5 => N18,
      O => OVtpg_inst_Row_10_GND_7_o_equal_8_o_10_1
    );
  OVtpg_inst_Row_10_GND_7_o_equal_5_o_10_1_SW0 : LUT3
    generic map(
      INIT => X"FD"
    )
    port map (
      I0 => OVtpg_inst_Row(3),
      I1 => OVtpg_inst_Row(5),
      I2 => OVtpg_inst_Row(4),
      O => N20
    );
  OVtpg_inst_Row_10_GND_7_o_equal_5_o_10_1 : LUT6
    generic map(
      INIT => X"0000000000000100"
    )
    port map (
      I0 => OVtpg_inst_Row(10),
      I1 => OVtpg_inst_Row(7),
      I2 => OVtpg_inst_Row(8),
      I3 => OVtpg_inst_Row(9),
      I4 => OVtpg_inst_Row(6),
      I5 => N20,
      O => OVtpg_inst_Row_10_GND_7_o_equal_5_o_10_1_96
    );
  OVtpg_inst_Mmux_pixel_out_12_pixel_out_23_mux_50_OUT3161 : LUT2
    generic map(
      INIT => X"8"
    )
    port map (
      I0 => OVtpg_inst_pmode(0),
      I1 => OVtpg_inst_n0133(0),
      O => OVtpg_inst_Mmux_pixel_out_12_pixel_out_23_mux_50_OUT3161_291
    );
  OVtpg_inst_Mmux_pixel_out_12_pixel_out_23_mux_50_OUT3163 : LUT6
    generic map(
      INIT => X"5555555554504400"
    )
    port map (
      I0 => OVtpg_inst_pmode(1),
      I1 => OVtpg_inst_Mmux_pixel_out_12_pixel_out_23_mux_50_OUT3111,
      I2 => OVtpg_inst_Mmux_pixel_out_12_pixel_out_23_mux_50_OUT3162_292,
      I3 => OVtpg_inst_Mmux_pixel_out_12_pixel_out_23_mux_50_OUT3161_291,
      I4 => OVtpg_inst_Mmux_pixel_out_12_pixel_out_23_mux_50_OUT3112,
      I5 => OVtpg_inst_Mmux_pixel_out_12_pixel_out_23_mux_50_OUT3113,
      O => OVtpg_inst_Mmux_pixel_out_12_pixel_out_23_mux_50_OUT3163_293
    );
  OVtpg_inst_Mmux_pixel_out_12_pixel_out_23_mux_50_OUT3167 : LUT6
    generic map(
      INIT => X"00000A00080EA0A0"
    )
    port map (
      I0 => OVtpg_inst_n0133(1),
      I1 => OVtpg_inst_n0133(2),
      I2 => OVtpg_inst_n0134(2),
      I3 => OVtpg_inst_n0133(0),
      I4 => OVtpg_inst_n0134(1),
      I5 => OVtpg_inst_n0134(0),
      O => OVtpg_inst_Mmux_pixel_out_12_pixel_out_23_mux_50_OUT3167_297
    );
  OVtpg_inst_Hsynci : FDR
    port map (
      C => clk_in_100,
      D => OVtpg_inst_Hsynci_glue_set_299,
      R => OVtpg_inst_n0262_200,
      Q => OVtpg_inst_Hsynci_234
    );
  OVtpg_inst_Active : FDR
    port map (
      C => clk_in_100,
      D => OVtpg_inst_Active_glue_set_300,
      R => OVtpg_inst_n0254_199,
      Q => OVtpg_inst_Active_235
    );
  OVtpg_inst_Hrefi : FDR
    port map (
      C => clk_in_100,
      D => OVtpg_inst_Hrefi_glue_set_301,
      R => OVtpg_inst_n0244_198,
      Q => OVtpg_inst_Hrefi_236
    );
  OVtpg_inst_Vsynci : FDR
    port map (
      C => clk_in_100,
      D => OVtpg_inst_Vsynci_glue_set,
      R => MRST,
      Q => OVtpg_inst_Vsynci_237
    );
  SIF_inst_vid_active_video : FDR
    port map (
      C => clk_in_50,
      D => SIF_inst_vid_active_video_glue_set_303,
      R => MRST,
      Q => NlwRenamedSig_OI_SIF_inst_vid_active_video
    );
  OVtpg_inst_Mcount_Col_cy_9_rt : LUT1
    generic map(
      INIT => X"2"
    )
    port map (
      I0 => OVtpg_inst_Col(9),
      O => OVtpg_inst_Mcount_Col_cy_9_rt_304
    );
  OVtpg_inst_Mcount_Col_cy_8_rt : LUT1
    generic map(
      INIT => X"2"
    )
    port map (
      I0 => OVtpg_inst_Col(8),
      O => OVtpg_inst_Mcount_Col_cy_8_rt_305
    );
  OVtpg_inst_Mcount_Col_cy_7_rt : LUT1
    generic map(
      INIT => X"2"
    )
    port map (
      I0 => OVtpg_inst_Col(7),
      O => OVtpg_inst_Mcount_Col_cy_7_rt_306
    );
  OVtpg_inst_Mcount_Col_cy_6_rt : LUT1
    generic map(
      INIT => X"2"
    )
    port map (
      I0 => OVtpg_inst_Col(6),
      O => OVtpg_inst_Mcount_Col_cy_6_rt_307
    );
  OVtpg_inst_Mcount_Col_cy_5_rt : LUT1
    generic map(
      INIT => X"2"
    )
    port map (
      I0 => OVtpg_inst_Col(5),
      O => OVtpg_inst_Mcount_Col_cy_5_rt_308
    );
  OVtpg_inst_Mcount_Col_cy_4_rt : LUT1
    generic map(
      INIT => X"2"
    )
    port map (
      I0 => OVtpg_inst_Col(4),
      O => OVtpg_inst_Mcount_Col_cy_4_rt_309
    );
  OVtpg_inst_Mcount_Col_cy_3_rt : LUT1
    generic map(
      INIT => X"2"
    )
    port map (
      I0 => OVtpg_inst_Col(3),
      O => OVtpg_inst_Mcount_Col_cy_3_rt_310
    );
  OVtpg_inst_Mcount_Col_cy_2_rt : LUT1
    generic map(
      INIT => X"2"
    )
    port map (
      I0 => OVtpg_inst_Col(2),
      O => OVtpg_inst_Mcount_Col_cy_2_rt_311
    );
  OVtpg_inst_Mcount_Col_cy_1_rt : LUT1
    generic map(
      INIT => X"2"
    )
    port map (
      I0 => OVtpg_inst_Col(1),
      O => OVtpg_inst_Mcount_Col_cy_1_rt_312
    );
  OVtpg_inst_Mcount_Row_cy_9_rt : LUT1
    generic map(
      INIT => X"2"
    )
    port map (
      I0 => OVtpg_inst_Row(9),
      O => OVtpg_inst_Mcount_Row_cy_9_rt_313
    );
  OVtpg_inst_Mcount_Row_cy_8_rt : LUT1
    generic map(
      INIT => X"2"
    )
    port map (
      I0 => OVtpg_inst_Row(8),
      O => OVtpg_inst_Mcount_Row_cy_8_rt_314
    );
  OVtpg_inst_Mcount_Row_cy_7_rt : LUT1
    generic map(
      INIT => X"2"
    )
    port map (
      I0 => OVtpg_inst_Row(7),
      O => OVtpg_inst_Mcount_Row_cy_7_rt_315
    );
  OVtpg_inst_Mcount_Row_cy_6_rt : LUT1
    generic map(
      INIT => X"2"
    )
    port map (
      I0 => OVtpg_inst_Row(6),
      O => OVtpg_inst_Mcount_Row_cy_6_rt_316
    );
  OVtpg_inst_Mcount_Row_cy_5_rt : LUT1
    generic map(
      INIT => X"2"
    )
    port map (
      I0 => OVtpg_inst_Row(5),
      O => OVtpg_inst_Mcount_Row_cy_5_rt_317
    );
  OVtpg_inst_Mcount_Row_cy_4_rt : LUT1
    generic map(
      INIT => X"2"
    )
    port map (
      I0 => OVtpg_inst_Row(4),
      O => OVtpg_inst_Mcount_Row_cy_4_rt_318
    );
  OVtpg_inst_Mcount_Row_cy_3_rt : LUT1
    generic map(
      INIT => X"2"
    )
    port map (
      I0 => OVtpg_inst_Row(3),
      O => OVtpg_inst_Mcount_Row_cy_3_rt_319
    );
  OVtpg_inst_Mcount_Row_cy_2_rt : LUT1
    generic map(
      INIT => X"2"
    )
    port map (
      I0 => OVtpg_inst_Row(2),
      O => OVtpg_inst_Mcount_Row_cy_2_rt_320
    );
  OVtpg_inst_Mcount_Row_cy_1_rt : LUT1
    generic map(
      INIT => X"2"
    )
    port map (
      I0 => OVtpg_inst_Row(1),
      O => OVtpg_inst_Mcount_Row_cy_1_rt_321
    );
  OVtpg_inst_Mcount_addr_cy_15_rt : LUT1
    generic map(
      INIT => X"2"
    )
    port map (
      I0 => NlwRenamedSig_OI_OVtpg_inst_addr(15),
      O => OVtpg_inst_Mcount_addr_cy_15_rt_322
    );
  OVtpg_inst_Mcount_addr_cy_14_rt : LUT1
    generic map(
      INIT => X"2"
    )
    port map (
      I0 => NlwRenamedSig_OI_OVtpg_inst_addr(14),
      O => OVtpg_inst_Mcount_addr_cy_14_rt_323
    );
  OVtpg_inst_Mcount_addr_cy_13_rt : LUT1
    generic map(
      INIT => X"2"
    )
    port map (
      I0 => NlwRenamedSig_OI_OVtpg_inst_addr(13),
      O => OVtpg_inst_Mcount_addr_cy_13_rt_324
    );
  OVtpg_inst_Mcount_addr_cy_12_rt : LUT1
    generic map(
      INIT => X"2"
    )
    port map (
      I0 => NlwRenamedSig_OI_OVtpg_inst_addr(12),
      O => OVtpg_inst_Mcount_addr_cy_12_rt_325
    );
  OVtpg_inst_Mcount_addr_cy_11_rt : LUT1
    generic map(
      INIT => X"2"
    )
    port map (
      I0 => NlwRenamedSig_OI_OVtpg_inst_addr(11),
      O => OVtpg_inst_Mcount_addr_cy_11_rt_326
    );
  OVtpg_inst_Mcount_addr_cy_10_rt : LUT1
    generic map(
      INIT => X"2"
    )
    port map (
      I0 => NlwRenamedSig_OI_OVtpg_inst_addr(10),
      O => OVtpg_inst_Mcount_addr_cy_10_rt_327
    );
  OVtpg_inst_Mcount_addr_cy_9_rt : LUT1
    generic map(
      INIT => X"2"
    )
    port map (
      I0 => NlwRenamedSig_OI_OVtpg_inst_addr(9),
      O => OVtpg_inst_Mcount_addr_cy_9_rt_328
    );
  OVtpg_inst_Mcount_addr_cy_8_rt : LUT1
    generic map(
      INIT => X"2"
    )
    port map (
      I0 => NlwRenamedSig_OI_OVtpg_inst_addr(8),
      O => OVtpg_inst_Mcount_addr_cy_8_rt_329
    );
  OVtpg_inst_Mcount_addr_cy_7_rt : LUT1
    generic map(
      INIT => X"2"
    )
    port map (
      I0 => NlwRenamedSig_OI_OVtpg_inst_addr(7),
      O => OVtpg_inst_Mcount_addr_cy_7_rt_330
    );
  OVtpg_inst_Mcount_addr_cy_6_rt : LUT1
    generic map(
      INIT => X"2"
    )
    port map (
      I0 => NlwRenamedSig_OI_OVtpg_inst_addr(6),
      O => OVtpg_inst_Mcount_addr_cy_6_rt_331
    );
  OVtpg_inst_Mcount_addr_cy_5_rt : LUT1
    generic map(
      INIT => X"2"
    )
    port map (
      I0 => NlwRenamedSig_OI_OVtpg_inst_addr(5),
      O => OVtpg_inst_Mcount_addr_cy_5_rt_332
    );
  OVtpg_inst_Mcount_addr_cy_4_rt : LUT1
    generic map(
      INIT => X"2"
    )
    port map (
      I0 => NlwRenamedSig_OI_OVtpg_inst_addr(4),
      O => OVtpg_inst_Mcount_addr_cy_4_rt_333
    );
  OVtpg_inst_Mcount_addr_cy_3_rt : LUT1
    generic map(
      INIT => X"2"
    )
    port map (
      I0 => NlwRenamedSig_OI_OVtpg_inst_addr(3),
      O => OVtpg_inst_Mcount_addr_cy_3_rt_334
    );
  OVtpg_inst_Mcount_addr_cy_2_rt : LUT1
    generic map(
      INIT => X"2"
    )
    port map (
      I0 => NlwRenamedSig_OI_OVtpg_inst_addr(2),
      O => OVtpg_inst_Mcount_addr_cy_2_rt_335
    );
  OVtpg_inst_Mcount_addr_cy_1_rt : LUT1
    generic map(
      INIT => X"2"
    )
    port map (
      I0 => NlwRenamedSig_OI_OVtpg_inst_addr(1),
      O => OVtpg_inst_Mcount_addr_cy_1_rt_336
    );
  OVtpg_inst_Mcount_Col_xor_10_rt : LUT1
    generic map(
      INIT => X"2"
    )
    port map (
      I0 => OVtpg_inst_Col(10),
      O => OVtpg_inst_Mcount_Col_xor_10_rt_337
    );
  OVtpg_inst_Mcount_Row_xor_10_rt : LUT1
    generic map(
      INIT => X"2"
    )
    port map (
      I0 => OVtpg_inst_Row(10),
      O => OVtpg_inst_Mcount_Row_xor_10_rt_338
    );
  OVtpg_inst_Mmux_pixel_out_12_pixel_out_23_mux_50_OUT3166 : LUT6
    generic map(
      INIT => X"FCCEA88ACEEC8AA8"
    )
    port map (
      I0 => OVtpg_inst_n0133(3),
      I1 => OVtpg_inst_n0134(3),
      I2 => OVtpg_inst_n0134(2),
      I3 => OVtpg_inst_n0134(1),
      I4 => OVtpg_inst_Mmux_pixel_out_12_pixel_out_23_mux_50_OUT3165_295,
      I5 => OVtpg_inst_n0134(0),
      O => OVtpg_inst_Mmux_pixel_out_12_pixel_out_23_mux_50_OUT3166_296
    );
  OVtpg_inst_Mmux_pixel_out_12_pixel_out_23_mux_50_OUT31131 : LUT4
    generic map(
      INIT => X"8880"
    )
    port map (
      I0 => OVtpg_inst_pmode(0),
      I1 => OVtpg_inst_n0133(3),
      I2 => OVtpg_inst_n0134(3),
      I3 => OVtpg_inst_n0134(2),
      O => OVtpg_inst_Mmux_pixel_out_12_pixel_out_23_mux_50_OUT3113
    );
  OVtpg_inst_Mmux_pixel_out_12_pixel_out_23_mux_50_OUT121_SW0 : LUT3
    generic map(
      INIT => X"80"
    )
    port map (
      I0 => OVtpg_inst_pmode(1),
      I1 => OVtpg_inst_pmode(0),
      I2 => N10,
      O => N32
    );
  OVtpg_inst_Mmux_pixel_out_12_pixel_out_23_mux_50_OUT121_SW1 : LUT5
    generic map(
      INIT => X"EAC0AA00"
    )
    port map (
      I0 => test_data(0),
      I1 => OVtpg_inst_pmode(1),
      I2 => OVtpg_inst_pmode(0),
      I3 => OVtpg_inst_Mmux_pixel_out_12_pixel_out_23_mux_50_OUT15,
      I4 => N10,
      O => N33
    );
  OVtpg_inst_Mmux_pixel_out_12_pixel_out_23_mux_50_OUT2 : LUT6
    generic map(
      INIT => X"FDFDFCFCFDB9FCB8"
    )
    port map (
      I0 => OVtpg_inst_pmode(2),
      I1 => OVtpg_inst_ClkDiv(1),
      I2 => N32,
      I3 => N33,
      I4 => OVtpg_inst_Mmux_pixel_out_12_pixel_out_23_mux_50_OUT317,
      I5 => OVtpg_inst_Mmux_pixel_out_12_pixel_out_23_mux_50_OUT316,
      O => OVtpg_inst_pixel_out_12_pixel_out_23_mux_50_OUT_1_Q
    );
  OVtpg_inst_Mmux_pixel_out_12_pixel_out_23_mux_50_OUT121_SW2 : LUT3
    generic map(
      INIT => X"80"
    )
    port map (
      I0 => OVtpg_inst_pmode(1),
      I1 => OVtpg_inst_pmode(0),
      I2 => N16,
      O => N35
    );
  OVtpg_inst_Mmux_pixel_out_12_pixel_out_23_mux_50_OUT121_SW3 : LUT5
    generic map(
      INIT => X"EAC0AA00"
    )
    port map (
      I0 => test_data(0),
      I1 => OVtpg_inst_pmode(1),
      I2 => OVtpg_inst_pmode(0),
      I3 => OVtpg_inst_Mmux_pixel_out_12_pixel_out_23_mux_50_OUT15,
      I4 => N16,
      O => N36
    );
  OVtpg_inst_Mmux_pixel_out_12_pixel_out_23_mux_50_OUT1 : LUT6
    generic map(
      INIT => X"FDFDFCFCFDB9FCB8"
    )
    port map (
      I0 => OVtpg_inst_pmode(2),
      I1 => OVtpg_inst_ClkDiv(1),
      I2 => N35,
      I3 => N36,
      I4 => OVtpg_inst_Mmux_pixel_out_12_pixel_out_23_mux_50_OUT317,
      I5 => OVtpg_inst_Mmux_pixel_out_12_pixel_out_23_mux_50_OUT316,
      O => OVtpg_inst_pixel_out_12_pixel_out_23_mux_50_OUT_0_Q
    );
  OVtpg_inst_Mmux_pixel_out_12_pixel_out_23_mux_50_OUT411_SW1 : LUT3
    generic map(
      INIT => X"F7"
    )
    port map (
      I0 => OVtpg_inst_pmode(1),
      I1 => OVtpg_inst_pmode(0),
      I2 => N12,
      O => N39
    );
  OVtpg_inst_Mmux_pixel_out_12_pixel_out_23_mux_50_OUT411_SW3 : LUT3
    generic map(
      INIT => X"F7"
    )
    port map (
      I0 => OVtpg_inst_pmode(1),
      I1 => OVtpg_inst_pmode(0),
      I2 => N14,
      O => N42
    );
  OVtpg_inst_Row_10_PWR_7_o_div_45_o_2_11 : LUT6
    generic map(
      INIT => X"F2F0F0F0F8F0F0F0"
    )
    port map (
      I0 => OVtpg_inst_Row(4),
      I1 => OVtpg_inst_Row(5),
      I2 => OVtpg_inst_Row_10_PWR_7_o_div_45_n0441_8_Q,
      I3 => OVtpg_inst_Row_10_PWR_7_o_div_45_Madd_a_10_GND_9_o_add_19_OUT_10_0_lut_7_Q,
      I4 => OVtpg_inst_Row_10_PWR_7_o_div_45_Madd_a_10_GND_9_o_add_19_OUT_10_0_lut_6_Q,
      I5 => OVtpg_inst_n0134(3),
      O => OVtpg_inst_n0134(2)
    );
  OVtpg_inst_Mmux_pixel_out_12_pixel_out_23_mux_50_OUT31612_SW0 : LUT6
    generic map(
      INIT => X"0C3BCCBBBBFEB3F2"
    )
    port map (
      I0 => OVtpg_inst_n0133(2),
      I1 => OVtpg_inst_n0134(2),
      I2 => OVtpg_inst_n0133(0),
      I3 => OVtpg_inst_n0134(1),
      I4 => N22,
      I5 => OVtpg_inst_n0134(0),
      O => N44
    );
  OVtpg_inst_Mmux_pixel_out_12_pixel_out_23_mux_50_OUT31111 : LUT6
    generic map(
      INIT => X"FFFFFFFFF8F0F0F0"
    )
    port map (
      I0 => OVtpg_inst_Row(4),
      I1 => OVtpg_inst_Row(5),
      I2 => OVtpg_inst_Row_10_PWR_7_o_div_45_n0441_8_Q,
      I3 => OVtpg_inst_Row_10_PWR_7_o_div_45_Madd_a_10_GND_9_o_add_19_OUT_10_0_lut_7_Q,
      I4 => OVtpg_inst_Row_10_PWR_7_o_div_45_Madd_a_10_GND_9_o_add_19_OUT_10_0_lut_6_Q,
      I5 => OVtpg_inst_n0134(3),
      O => OVtpg_inst_Mmux_pixel_out_12_pixel_out_23_mux_50_OUT3111
    );
  OVtpg_inst_Row_10_PWR_7_o_div_45_Mmux_n044181 : LUT6
    generic map(
      INIT => X"9886966696669666"
    )
    port map (
      I0 => OVtpg_inst_Row(10),
      I1 => OVtpg_inst_Row(6),
      I2 => OVtpg_inst_Row(9),
      I3 => OVtpg_inst_Row(5),
      I4 => OVtpg_inst_Row(8),
      I5 => OVtpg_inst_Row(7),
      O => OVtpg_inst_Row_10_PWR_7_o_div_45_Madd_a_10_GND_9_o_add_19_OUT_10_0_lut_6_Q
    );
  OVtpg_inst_Row_10_PWR_7_o_div_45_o_0_121 : LUT5
    generic map(
      INIT => X"79999999"
    )
    port map (
      I0 => OVtpg_inst_Row(6),
      I1 => OVtpg_inst_Row(10),
      I2 => OVtpg_inst_Row(7),
      I3 => OVtpg_inst_Row(8),
      I4 => OVtpg_inst_Row(9),
      O => OVtpg_inst_Row_10_PWR_7_o_div_45_o_0_12
    );
  OVtpg_inst_Mmux_pixel_out_12_pixel_out_23_mux_50_OUT83 : LUT6
    generic map(
      INIT => X"FFDDFBD9FFCCFBC8"
    )
    port map (
      I0 => OVtpg_inst_pmode(2),
      I1 => OVtpg_inst_ClkDiv(1),
      I2 => N49,
      I3 => N48,
      I4 => OVtpg_inst_Mmux_pixel_out_12_pixel_out_23_mux_50_OUT317,
      I5 => OVtpg_inst_Mmux_pixel_out_12_pixel_out_23_mux_50_OUT4112,
      O => OVtpg_inst_pixel_out_12_pixel_out_23_mux_50_OUT_7_Q
    );
  OVtpg_inst_Row_10_PWR_7_o_div_45_o_1_11_SW0 : LUT2
    generic map(
      INIT => X"8"
    )
    port map (
      I0 => OVtpg_inst_Row(3),
      I1 => OVtpg_inst_Row_10_PWR_7_o_div_45_o_0_11,
      O => N55
    );
  OVtpg_inst_Row_10_PWR_7_o_div_45_o_1_12 : LUT6
    generic map(
      INIT => X"AEFEEA6AAAFAAA2A"
    )
    port map (
      I0 => OVtpg_inst_Row_10_PWR_7_o_div_45_Madd_a_10_GND_9_o_add_19_OUT_10_0_lut_7_Q,
      I1 => OVtpg_inst_Row_10_PWR_7_o_div_45_Madd_a_10_GND_9_o_add_19_OUT_10_0_lut_6_Q,
      I2 => OVtpg_inst_Row(4),
      I3 => N56,
      I4 => OVtpg_inst_Row_10_PWR_7_o_div_45_n0441_8_Q,
      I5 => N55,
      O => OVtpg_inst_n0134(1)
    );
  OVtpg_inst_Row_10_PWR_7_o_div_45_o_0_111 : LUT6
    generic map(
      INIT => X"9886666666666666"
    )
    port map (
      I0 => OVtpg_inst_Row(5),
      I1 => OVtpg_inst_Row(9),
      I2 => OVtpg_inst_Row(6),
      I3 => OVtpg_inst_Row(10),
      I4 => OVtpg_inst_Row(7),
      I5 => OVtpg_inst_Row(8),
      O => OVtpg_inst_Row_10_PWR_7_o_div_45_o_0_11
    );
  OVtpg_inst_Mmux_pixel_out_12_pixel_out_23_mux_50_OUT3165 : LUT3
    generic map(
      INIT => X"96"
    )
    port map (
      I0 => OVtpg_inst_n0133(1),
      I1 => OVtpg_inst_n0133(2),
      I2 => OVtpg_inst_n0133(0),
      O => OVtpg_inst_Mmux_pixel_out_12_pixel_out_23_mux_50_OUT3165_295
    );
  OVtpg_inst_Col_10_PWR_7_o_div_44_o_1_1 : LUT6
    generic map(
      INIT => X"03E880FEFE033F80"
    )
    port map (
      I0 => OVtpg_inst_Col(5),
      I1 => OVtpg_inst_Col(6),
      I2 => OVtpg_inst_Col(10),
      I3 => OVtpg_inst_Col(9),
      I4 => OVtpg_inst_Col(8),
      I5 => OVtpg_inst_Col(7),
      O => OVtpg_inst_n0133(1)
    );
  OVtpg_inst_Row_10_PWR_7_o_div_45_Mmux_n044192 : LUT6
    generic map(
      INIT => X"554646AA552A2AAA"
    )
    port map (
      I0 => OVtpg_inst_Row(7),
      I1 => OVtpg_inst_Row(5),
      I2 => OVtpg_inst_Row(8),
      I3 => OVtpg_inst_Row(10),
      I4 => OVtpg_inst_Row(6),
      I5 => OVtpg_inst_Row(9),
      O => OVtpg_inst_Row_10_PWR_7_o_div_45_Madd_a_10_GND_9_o_add_19_OUT_10_0_lut_7_Q
    );
  OVtpg_inst_Row_10_PWR_7_o_div_45_Mmux_n0441101 : LUT6
    generic map(
      INIT => X"554242AAAAAAAAAA"
    )
    port map (
      I0 => OVtpg_inst_Row(8),
      I1 => OVtpg_inst_Row(9),
      I2 => OVtpg_inst_Row(5),
      I3 => OVtpg_inst_Row(10),
      I4 => OVtpg_inst_Row(6),
      I5 => OVtpg_inst_Row(7),
      O => OVtpg_inst_Row_10_PWR_7_o_div_45_n0441_8_Q
    );
  OVtpg_inst_Mmux_pixel_out_12_pixel_out_23_mux_50_OUT31613_SW0 : LUT5
    generic map(
      INIT => X"CCFFCCFE"
    )
    port map (
      I0 => OVtpg_inst_n0133(3),
      I1 => OVtpg_inst_n0134(3),
      I2 => OVtpg_inst_n0133(1),
      I3 => OVtpg_inst_Mmux_pixel_out_12_pixel_out_23_mux_50_OUT3167_297,
      I4 => N44,
      O => N91
    );
  OVtpg_inst_Mmux_pixel_out_12_pixel_out_23_mux_50_OUT31613 : LUT6
    generic map(
      INIT => X"FFA0FFA8FFA2FFAA"
    )
    port map (
      I0 => OVtpg_inst_Mmux_pixel_out_12_pixel_out_23_mux_50_OUT3164,
      I1 => OVtpg_inst_Mmux_pixel_out_12_pixel_out_23_mux_50_OUT3169_298,
      I2 => OVtpg_inst_Mmux_pixel_out_12_pixel_out_23_mux_50_OUT3166_296,
      I3 => OVtpg_inst_Mmux_pixel_out_12_pixel_out_23_mux_50_OUT3163_293,
      I4 => N92,
      I5 => N91,
      O => OVtpg_inst_Mmux_pixel_out_12_pixel_out_23_mux_50_OUT316
    );
  OVtpg_inst_Mmux_pixel_out_12_pixel_out_23_mux_50_OUT41128_SW0 : LUT5
    generic map(
      INIT => X"FDDCEF0A"
    )
    port map (
      I0 => OVtpg_inst_n0133(2),
      I1 => OVtpg_inst_n0134(3),
      I2 => OVtpg_inst_n0133(1),
      I3 => OVtpg_inst_n0133(0),
      I4 => OVtpg_inst_n0134(2),
      O => N94
    );
  OVtpg_inst_Mmux_pixel_out_12_pixel_out_23_mux_50_OUT41128_SW1 : LUT4
    generic map(
      INIT => X"FCEA"
    )
    port map (
      I0 => OVtpg_inst_n0133(2),
      I1 => OVtpg_inst_n0134(3),
      I2 => OVtpg_inst_n0133(0),
      I3 => OVtpg_inst_n0134(2),
      O => N95
    );
  OVtpg_inst_Mmux_pixel_out_12_pixel_out_23_mux_50_OUT41128 : LUT5
    generic map(
      INIT => X"00401050"
    )
    port map (
      I0 => OVtpg_inst_n0133(3),
      I1 => OVtpg_inst_n0134(1),
      I2 => OVtpg_inst_n0134(0),
      I3 => N95,
      I4 => N94,
      O => OVtpg_inst_Mmux_pixel_out_12_pixel_out_23_mux_50_OUT41128_271
    );
  OVtpg_inst_Mmux_pixel_out_12_pixel_out_23_mux_50_OUT41126_SW0 : LUT4
    generic map(
      INIT => X"1105"
    )
    port map (
      I0 => OVtpg_inst_n0133(3),
      I1 => OVtpg_inst_n0133(2),
      I2 => OVtpg_inst_n0133(0),
      I3 => OVtpg_inst_n0134(2),
      O => N97
    );
  OVtpg_inst_Mmux_pixel_out_12_pixel_out_23_mux_50_OUT41126_SW1 : LUT5
    generic map(
      INIT => X"10510445"
    )
    port map (
      I0 => OVtpg_inst_n0133(3),
      I1 => OVtpg_inst_n0133(2),
      I2 => OVtpg_inst_n0133(1),
      I3 => OVtpg_inst_n0133(0),
      I4 => OVtpg_inst_n0134(2),
      O => N98
    );
  OVtpg_inst_Mmux_pixel_out_12_pixel_out_23_mux_50_OUT41126 : LUT6
    generic map(
      INIT => X"F0F0F0F4F0F1F0F5"
    )
    port map (
      I0 => OVtpg_inst_n0134(3),
      I1 => OVtpg_inst_n0134(1),
      I2 => OVtpg_inst_Mmux_pixel_out_12_pixel_out_23_mux_50_OUT41124_269,
      I3 => OVtpg_inst_n0134(0),
      I4 => N98,
      I5 => N97,
      O => OVtpg_inst_Mmux_pixel_out_12_pixel_out_23_mux_50_OUT41126_270
    );
  OVtpg_inst_Row_10_PWR_7_o_div_45_o_1_11_SW1 : LUT6
    generic map(
      INIT => X"7FFFF99FF99FF99F"
    )
    port map (
      I0 => OVtpg_inst_Row(9),
      I1 => OVtpg_inst_Row(5),
      I2 => OVtpg_inst_Row(6),
      I3 => OVtpg_inst_Row(10),
      I4 => OVtpg_inst_Row(7),
      I5 => OVtpg_inst_Row(8),
      O => N56
    );
  OVtpg_inst_Mmux_pixel_out_12_pixel_out_23_mux_50_OUT3177_SW2 : LUT4
    generic map(
      INIT => X"FA11"
    )
    port map (
      I0 => OVtpg_inst_n0133(3),
      I1 => OVtpg_inst_n0133(2),
      I2 => OVtpg_inst_n0133(0),
      I3 => OVtpg_inst_n0134(2),
      O => N100
    );
  OVtpg_inst_Mmux_pixel_out_12_pixel_out_23_mux_50_OUT3177_SW3 : LUT5
    generic map(
      INIT => X"EFAE0445"
    )
    port map (
      I0 => OVtpg_inst_n0133(3),
      I1 => OVtpg_inst_n0133(2),
      I2 => OVtpg_inst_n0133(1),
      I3 => OVtpg_inst_n0133(0),
      I4 => OVtpg_inst_n0134(2),
      O => N101
    );
  OVtpg_inst_Mmux_pixel_out_12_pixel_out_23_mux_50_OUT3177_SW4 : LUT5
    generic map(
      INIT => X"0445EFAE"
    )
    port map (
      I0 => OVtpg_inst_n0133(3),
      I1 => OVtpg_inst_n0133(2),
      I2 => OVtpg_inst_n0133(1),
      I3 => OVtpg_inst_n0133(0),
      I4 => OVtpg_inst_n0134(2),
      O => N102
    );
  OVtpg_inst_Mmux_pixel_out_12_pixel_out_23_mux_50_OUT3177 : LUT6
    generic map(
      INIT => X"5140D9C87362FBEA"
    )
    port map (
      I0 => OVtpg_inst_n0134(1),
      I1 => OVtpg_inst_n0134(0),
      I2 => N101,
      I3 => N100,
      I4 => N103,
      I5 => N102,
      O => OVtpg_inst_Mmux_pixel_out_12_pixel_out_23_mux_50_OUT3177_264
    );
  OVtpg_inst_Mmux_pixel_out_12_pixel_out_23_mux_50_OUT3167_SW0 : LUT4
    generic map(
      INIT => X"CEEE"
    )
    port map (
      I0 => OVtpg_inst_n0133(3),
      I1 => OVtpg_inst_n0134(3),
      I2 => OVtpg_inst_n0133(1),
      I3 => OVtpg_inst_n0134(2),
      O => N105
    );
  OVtpg_inst_Mmux_pixel_out_12_pixel_out_23_mux_50_OUT3167_SW1 : LUT5
    generic map(
      INIT => X"EEEECEEE"
    )
    port map (
      I0 => OVtpg_inst_n0133(3),
      I1 => OVtpg_inst_n0134(3),
      I2 => OVtpg_inst_n0133(1),
      I3 => OVtpg_inst_n0133(0),
      I4 => OVtpg_inst_n0134(2),
      O => N106
    );
  OVtpg_inst_Mmux_pixel_out_12_pixel_out_23_mux_50_OUT3167_SW2 : LUT6
    generic map(
      INIT => X"FAFAFAFAF2FAF0F2"
    )
    port map (
      I0 => OVtpg_inst_n0133(3),
      I1 => OVtpg_inst_n0133(2),
      I2 => OVtpg_inst_n0134(3),
      I3 => OVtpg_inst_n0133(1),
      I4 => OVtpg_inst_n0133(0),
      I5 => OVtpg_inst_n0134(2),
      O => N107
    );
  OVtpg_inst_Mmux_pixel_out_12_pixel_out_23_mux_50_OUT31613_SW1 : LUT6
    generic map(
      INIT => X"BFBC8F8CB3B08380"
    )
    port map (
      I0 => N108,
      I1 => OVtpg_inst_n0134(1),
      I2 => OVtpg_inst_n0134(0),
      I3 => N105,
      I4 => N106,
      I5 => N107,
      O => N92
    );
  OVtpg_inst_Mmux_pixel_out_12_pixel_out_23_mux_50_OUT5 : LUT6
    generic map(
      INIT => X"55115F1BF5B1FFBB"
    )
    port map (
      I0 => OVtpg_inst_ClkDiv(1),
      I1 => N110,
      I2 => N91,
      I3 => OVtpg_inst_Mmux_pixel_out_12_pixel_out_23_mux_50_OUT4112,
      I4 => N111,
      I5 => N112,
      O => OVtpg_inst_pixel_out_12_pixel_out_23_mux_50_OUT_4_Q
    );
  OVtpg_inst_Mmux_pixel_out_12_pixel_out_23_mux_50_OUT4 : LUT6
    generic map(
      INIT => X"55115F1BF5B1FFBB"
    )
    port map (
      I0 => OVtpg_inst_ClkDiv(1),
      I1 => N114,
      I2 => N91,
      I3 => OVtpg_inst_Mmux_pixel_out_12_pixel_out_23_mux_50_OUT4112,
      I4 => N115,
      I5 => N116,
      O => OVtpg_inst_pixel_out_12_pixel_out_23_mux_50_OUT_3_Q
    );
  OVtpg_inst_Mmux_pixel_out_12_pixel_out_23_mux_50_OUT3162 : LUT5
    generic map(
      INIT => X"00003B9D"
    )
    port map (
      I0 => OVtpg_inst_Col(10),
      I1 => OVtpg_inst_Col(9),
      I2 => OVtpg_inst_Col(7),
      I3 => OVtpg_inst_Col(8),
      I4 => OVtpg_inst_n0133(0),
      O => OVtpg_inst_Mmux_pixel_out_12_pixel_out_23_mux_50_OUT3162_292
    );
  OVtpg_inst_Mmux_pixel_out_12_pixel_out_23_mux_50_OUT73 : LUT6
    generic map(
      INIT => X"FFFFFFB3FFCCFF80"
    )
    port map (
      I0 => test_data(4),
      I1 => OVtpg_inst_ClkDiv(1),
      I2 => OVtpg_inst_Mmux_pixel_out_12_pixel_out_23_mux_50_OUT15,
      I3 => OVtpg_inst_Mmux_pixel_out_12_pixel_out_23_mux_50_OUT71_277,
      I4 => OVtpg_inst_Mmux_pixel_out_12_pixel_out_23_mux_50_OUT317,
      I5 => OVtpg_inst_Mmux_pixel_out_12_pixel_out_23_mux_50_OUT4112,
      O => OVtpg_inst_pixel_out_12_pixel_out_23_mux_50_OUT_6_Q
    );
  OVtpg_inst_Mmux_pixel_out_12_pixel_out_23_mux_50_OUT63 : LUT6
    generic map(
      INIT => X"FFFFFFB3FFCCFF80"
    )
    port map (
      I0 => test_data(4),
      I1 => OVtpg_inst_ClkDiv(1),
      I2 => OVtpg_inst_Mmux_pixel_out_12_pixel_out_23_mux_50_OUT15,
      I3 => OVtpg_inst_Mmux_pixel_out_12_pixel_out_23_mux_50_OUT61_279,
      I4 => OVtpg_inst_Mmux_pixel_out_12_pixel_out_23_mux_50_OUT317,
      I5 => OVtpg_inst_Mmux_pixel_out_12_pixel_out_23_mux_50_OUT4112,
      O => OVtpg_inst_pixel_out_12_pixel_out_23_mux_50_OUT_5_Q
    );
  OVtpg_inst_Mmux_pixel_out_12_pixel_out_23_mux_50_OUT3169 : LUT6
    generic map(
      INIT => X"0000406805004068"
    )
    port map (
      I0 => OVtpg_inst_n0133(2),
      I1 => OVtpg_inst_n0133(1),
      I2 => OVtpg_inst_n0133(0),
      I3 => OVtpg_inst_n0134(2),
      I4 => OVtpg_inst_n0134(1),
      I5 => OVtpg_inst_n0134(0),
      O => OVtpg_inst_Mmux_pixel_out_12_pixel_out_23_mux_50_OUT3169_298
    );
  OVtpg_inst_Mmux_pixel_out_12_pixel_out_23_mux_50_OUT31613_SW2 : LUT6
    generic map(
      INIT => X"1111333301110333"
    )
    port map (
      I0 => test_data(8),
      I1 => OVtpg_inst_pmode(2),
      I2 => OVtpg_inst_pmode(1),
      I3 => OVtpg_inst_pmode(0),
      I4 => OVtpg_inst_Mmux_pixel_out_12_pixel_out_23_mux_50_OUT15,
      I5 => N12,
      O => N110
    );
  OVtpg_inst_Mmux_pixel_out_12_pixel_out_23_mux_50_OUT31613_SW5 : LUT6
    generic map(
      INIT => X"1111333301110333"
    )
    port map (
      I0 => test_data(8),
      I1 => OVtpg_inst_pmode(2),
      I2 => OVtpg_inst_pmode(1),
      I3 => OVtpg_inst_pmode(0),
      I4 => OVtpg_inst_Mmux_pixel_out_12_pixel_out_23_mux_50_OUT15,
      I5 => N14,
      O => N114
    );
  OVtpg_inst_Mmux_pixel_out_12_pixel_out_23_mux_50_OUT82111 : LUT6
    generic map(
      INIT => X"8888880888888888"
    )
    port map (
      I0 => OVtpg_inst_pmode(0),
      I1 => OVtpg_inst_pmode(1),
      I2 => OVtpg_inst_Inside1_287,
      I3 => OVtpg_inst_Col(9),
      I4 => OVtpg_inst_Col(10),
      I5 => OVtpg_inst_Inside2_288,
      O => OVtpg_inst_Mmux_pixel_out_12_pixel_out_23_mux_50_OUT15
    );
  OVtpg_inst_Mmux_pixel_out_12_pixel_out_23_mux_50_OUT41124 : LUT6
    generic map(
      INIT => X"0000000028A8222A"
    )
    port map (
      I0 => OVtpg_inst_n0134(3),
      I1 => OVtpg_inst_Col(9),
      I2 => OVtpg_inst_Col(8),
      I3 => OVtpg_inst_Col(7),
      I4 => OVtpg_inst_Col(10),
      I5 => OVtpg_inst_n0133(0),
      O => OVtpg_inst_Mmux_pixel_out_12_pixel_out_23_mux_50_OUT41124_269
    );
  OVtpg_inst_Mmux_pixel_out_12_pixel_out_23_mux_50_OUT3177_SW5 : LUT6
    generic map(
      INIT => X"FFFFFFFFFFFFC462"
    )
    port map (
      I0 => OVtpg_inst_Col(10),
      I1 => OVtpg_inst_Col(9),
      I2 => OVtpg_inst_Col(7),
      I3 => OVtpg_inst_Col(8),
      I4 => OVtpg_inst_n0133(0),
      I5 => OVtpg_inst_n0134(2),
      O => N103
    );
  OVtpg_inst_Mmux_pixel_out_12_pixel_out_23_mux_50_OUT31613_SW3 : MUXF7
    port map (
      I0 => N124,
      I1 => N125,
      S => OVtpg_inst_Mmux_pixel_out_12_pixel_out_23_mux_50_OUT3169_298,
      O => N111
    );
  OVtpg_inst_Mmux_pixel_out_12_pixel_out_23_mux_50_OUT31613_SW3_G : LUT6
    generic map(
      INIT => X"A0A0A0A0B0F0B0B0"
    )
    port map (
      I0 => OVtpg_inst_pmode(2),
      I1 => OVtpg_inst_Mmux_pixel_out_12_pixel_out_23_mux_50_OUT3164,
      I2 => N39,
      I3 => OVtpg_inst_Mmux_pixel_out_12_pixel_out_23_mux_50_OUT3166_296,
      I4 => N92,
      I5 => OVtpg_inst_Mmux_pixel_out_12_pixel_out_23_mux_50_OUT3163_293,
      O => N125
    );
  OVtpg_inst_Mmux_pixel_out_12_pixel_out_23_mux_50_OUT31613_SW4 : MUXF7
    port map (
      I0 => N126,
      I1 => N127,
      S => OVtpg_inst_Mmux_pixel_out_12_pixel_out_23_mux_50_OUT3169_298,
      O => N112
    );
  OVtpg_inst_Mmux_pixel_out_12_pixel_out_23_mux_50_OUT31613_SW4_G : LUT6
    generic map(
      INIT => X"A0A0A0A0B0F0B0B0"
    )
    port map (
      I0 => OVtpg_inst_pmode(2),
      I1 => OVtpg_inst_Mmux_pixel_out_12_pixel_out_23_mux_50_OUT3164,
      I2 => N39,
      I3 => OVtpg_inst_Mmux_pixel_out_12_pixel_out_23_mux_50_OUT3166_296,
      I4 => N92,
      I5 => OVtpg_inst_Mmux_pixel_out_12_pixel_out_23_mux_50_OUT3163_293,
      O => N127
    );
  OVtpg_inst_Mmux_pixel_out_12_pixel_out_23_mux_50_OUT31613_SW6 : MUXF7
    port map (
      I0 => N128,
      I1 => N129,
      S => OVtpg_inst_Mmux_pixel_out_12_pixel_out_23_mux_50_OUT3169_298,
      O => N115
    );
  OVtpg_inst_Mmux_pixel_out_12_pixel_out_23_mux_50_OUT31613_SW6_G : LUT6
    generic map(
      INIT => X"A0A0A0A0B0F0B0B0"
    )
    port map (
      I0 => OVtpg_inst_pmode(2),
      I1 => OVtpg_inst_Mmux_pixel_out_12_pixel_out_23_mux_50_OUT3164,
      I2 => N42,
      I3 => OVtpg_inst_Mmux_pixel_out_12_pixel_out_23_mux_50_OUT3166_296,
      I4 => N92,
      I5 => OVtpg_inst_Mmux_pixel_out_12_pixel_out_23_mux_50_OUT3163_293,
      O => N129
    );
  OVtpg_inst_Mmux_pixel_out_12_pixel_out_23_mux_50_OUT31613_SW7 : MUXF7
    port map (
      I0 => N130,
      I1 => N131,
      S => OVtpg_inst_Mmux_pixel_out_12_pixel_out_23_mux_50_OUT3169_298,
      O => N116
    );
  OVtpg_inst_Mmux_pixel_out_12_pixel_out_23_mux_50_OUT31613_SW7_G : LUT6
    generic map(
      INIT => X"A0A0A0A0B0F0B0B0"
    )
    port map (
      I0 => OVtpg_inst_pmode(2),
      I1 => OVtpg_inst_Mmux_pixel_out_12_pixel_out_23_mux_50_OUT3164,
      I2 => N42,
      I3 => OVtpg_inst_Mmux_pixel_out_12_pixel_out_23_mux_50_OUT3166_296,
      I4 => N92,
      I5 => OVtpg_inst_Mmux_pixel_out_12_pixel_out_23_mux_50_OUT3163_293,
      O => N131
    );
  OVtpg_inst_Hsynci_glue_set : LUT3
    generic map(
      INIT => X"FD"
    )
    port map (
      I0 => locked_in,
      I1 => OVtpg_inst_Hsynci_234,
      I2 => OVtpg_inst_n0358_inv_184,
      O => OVtpg_inst_Hsynci_glue_set_299
    );
  OVtpg_inst_Hrefi_glue_set : LUT6
    generic map(
      INIT => X"FBBBBBBBBBBBBBBB"
    )
    port map (
      I0 => OVtpg_inst_Hrefi_236,
      I1 => locked_in,
      I2 => OVtpg_inst_ClkDiv(0),
      I3 => OVtpg_inst_ClkDiv(1),
      I4 => OVtpg_inst_Col_10_GND_7_o_equal_4_o,
      I5 => OVtpg_inst_Active_235,
      O => OVtpg_inst_Hrefi_glue_set_301
    );
  OVtpg_inst_n0395_inv3_SW0 : LUT6
    generic map(
      INIT => X"FFBFFFFFFFFFFFFF"
    )
    port map (
      I0 => OVtpg_inst_Col(8),
      I1 => OVtpg_inst_Col(1),
      I2 => OVtpg_inst_Col(2),
      I3 => OVtpg_inst_Col(10),
      I4 => OVtpg_inst_Col(3),
      I5 => OVtpg_inst_Col(9),
      O => N132
    );
  OVtpg_inst_n0395_inv3 : LUT6
    generic map(
      INIT => X"FFFF9FFFFFFFFBFF"
    )
    port map (
      I0 => OVtpg_inst_Col(4),
      I1 => OVtpg_inst_Col(7),
      I2 => OVtpg_inst_Col(6),
      I3 => OVtpg_inst_Col(0),
      I4 => N132,
      I5 => OVtpg_inst_Col(5),
      O => OVtpg_inst_n0395_inv3_275
    );
  OVtpg_inst_n0254_SW1 : LUT4
    generic map(
      INIT => X"BFFF"
    )
    port map (
      I0 => OVtpg_inst_Row(5),
      I1 => OVtpg_inst_Row(2),
      I2 => OVtpg_inst_Row(4),
      I3 => locked_in,
      O => N134
    );
  OVtpg_inst_n0254 : LUT6
    generic map(
      INIT => X"2000000000000000"
    )
    port map (
      I0 => OVtpg_inst_ClkDiv(1),
      I1 => N134,
      I2 => OVtpg_inst_Col_10_GND_7_o_equal_4_o,
      I3 => OVtpg_inst_Row_10_GND_7_o_equal_8_o_10_1,
      I4 => OVtpg_inst_Row(1),
      I5 => OVtpg_inst_ClkDiv(0),
      O => OVtpg_inst_n0254_199
    );
  OVtpg_inst_Mmux_pixel_out_12_pixel_out_23_mux_50_OUT3171 : LUT6
    generic map(
      INIT => X"28202828A2822820"
    )
    port map (
      I0 => OVtpg_inst_pmode(0),
      I1 => OVtpg_inst_Col(8),
      I2 => OVtpg_inst_Col(10),
      I3 => OVtpg_inst_Col(6),
      I4 => OVtpg_inst_Col(9),
      I5 => OVtpg_inst_Col(7),
      O => OVtpg_inst_Mmux_pixel_out_12_pixel_out_23_mux_50_OUT3171_261
    );
  OVtpg_inst_Mcount_Col_val1 : LUT4
    generic map(
      INIT => X"D555"
    )
    port map (
      I0 => locked_in,
      I1 => OVtpg_inst_ClkDiv(0),
      I2 => OVtpg_inst_Col_10_GND_7_o_equal_4_o,
      I3 => OVtpg_inst_ClkDiv(1),
      O => OVtpg_inst_Mcount_Col_val
    );
  OVtpg_inst_n0262 : LUT5
    generic map(
      INIT => X"00000200"
    )
    port map (
      I0 => OVtpg_inst_Col_10_GND_7_o_equal_4_o_10_1,
      I1 => OVtpg_inst_Col(6),
      I2 => OVtpg_inst_Col(8),
      I3 => OVtpg_inst_Col(7),
      I4 => N6,
      O => OVtpg_inst_n0262_200
    );
  OVtpg_inst_Mmux_pixel_out_12_pixel_out_23_mux_50_OUT821_SW0 : LUT3
    generic map(
      INIT => X"80"
    )
    port map (
      I0 => OVtpg_inst_pmode(1),
      I1 => OVtpg_inst_pmode(0),
      I2 => OVtpg_inst_Mmux_pixel_out_12_pixel_out_23_mux_50_OUT8,
      O => N48
    );
  OVtpg_inst_Mmux_pixel_out_12_pixel_out_23_mux_50_OUT821_SW1 : LUT5
    generic map(
      INIT => X"F8888888"
    )
    port map (
      I0 => OVtpg_inst_Mmux_pixel_out_12_pixel_out_23_mux_50_OUT15,
      I1 => test_data(4),
      I2 => OVtpg_inst_pmode(0),
      I3 => OVtpg_inst_pmode(1),
      I4 => OVtpg_inst_Mmux_pixel_out_12_pixel_out_23_mux_50_OUT8,
      O => N49
    );
  OVtpg_inst_Mmux_pixel_out_12_pixel_out_23_mux_50_OUT3167_SW3 : LUT5
    generic map(
      INIT => X"FFFF91A8"
    )
    port map (
      I0 => OVtpg_inst_Col(9),
      I1 => OVtpg_inst_Col(8),
      I2 => OVtpg_inst_Col(7),
      I3 => OVtpg_inst_Col(10),
      I4 => OVtpg_inst_n0134(3),
      O => N108
    );
  SIF_inst_vid_active_video_glue_set : LUT3
    generic map(
      INIT => X"A8"
    )
    port map (
      I0 => OVtpg_inst_HREF_61,
      I1 => NlwRenamedSig_OI_SIF_inst_vid_active_video,
      I2 => SIF_inst_oddpix_252,
      O => SIF_inst_vid_active_video_glue_set_303
    );
  OVtpg_inst_Mmux_pixel_out_12_pixel_out_23_mux_50_OUT3172 : LUT5
    generic map(
      INIT => X"41414159"
    )
    port map (
      I0 => OVtpg_inst_Col(9),
      I1 => OVtpg_inst_Col(10),
      I2 => OVtpg_inst_Col(8),
      I3 => OVtpg_inst_Col(7),
      I4 => OVtpg_inst_Col(6),
      O => OVtpg_inst_Mmux_pixel_out_12_pixel_out_23_mux_50_OUT3172_262
    );
  OVtpg_inst_Mmux_pixel_out_12_pixel_out_23_mux_50_OUT41122 : LUT6
    generic map(
      INIT => X"0509158914815491"
    )
    port map (
      I0 => OVtpg_inst_Col(9),
      I1 => OVtpg_inst_Col(10),
      I2 => OVtpg_inst_Col(7),
      I3 => OVtpg_inst_Col(8),
      I4 => OVtpg_inst_Col(5),
      I5 => OVtpg_inst_Col(6),
      O => OVtpg_inst_Mmux_pixel_out_12_pixel_out_23_mux_50_OUT41122_267
    );
  OVtpg_inst_Mmux_pixel_out_12_pixel_out_23_mux_50_OUT3178 : LUT5
    generic map(
      INIT => X"FFFB6664"
    )
    port map (
      I0 => OVtpg_inst_Col(8),
      I1 => OVtpg_inst_Col(10),
      I2 => OVtpg_inst_Col(6),
      I3 => OVtpg_inst_Col(7),
      I4 => OVtpg_inst_Col(9),
      O => OVtpg_inst_Mmux_pixel_out_12_pixel_out_23_mux_50_OUT3178_265
    );
  OVtpg_inst_Mmux_pixel_out_12_pixel_out_23_mux_50_OUT31613_SW3_F : LUT5
    generic map(
      INIT => X"AA2AFB3B"
    )
    port map (
      I0 => OVtpg_inst_pmode(2),
      I1 => OVtpg_inst_pmode(1),
      I2 => OVtpg_inst_pmode(0),
      I3 => N12,
      I4 => OVtpg_inst_Mmux_pixel_out_12_pixel_out_23_mux_50_OUT3163_293,
      O => N124
    );
  OVtpg_inst_Mmux_pixel_out_12_pixel_out_23_mux_50_OUT31613_SW4_F : LUT6
    generic map(
      INIT => X"AA2AAA2AFB3BFF3F"
    )
    port map (
      I0 => OVtpg_inst_pmode(2),
      I1 => OVtpg_inst_pmode(1),
      I2 => OVtpg_inst_pmode(0),
      I3 => N12,
      I4 => OVtpg_inst_Mmux_pixel_out_12_pixel_out_23_mux_50_OUT3166_296,
      I5 => OVtpg_inst_Mmux_pixel_out_12_pixel_out_23_mux_50_OUT3163_293,
      O => N126
    );
  OVtpg_inst_Mmux_pixel_out_12_pixel_out_23_mux_50_OUT31613_SW6_F : LUT5
    generic map(
      INIT => X"AA2AFB3B"
    )
    port map (
      I0 => OVtpg_inst_pmode(2),
      I1 => OVtpg_inst_pmode(1),
      I2 => OVtpg_inst_pmode(0),
      I3 => N14,
      I4 => OVtpg_inst_Mmux_pixel_out_12_pixel_out_23_mux_50_OUT3163_293,
      O => N128
    );
  OVtpg_inst_Mmux_pixel_out_12_pixel_out_23_mux_50_OUT31613_SW7_F : LUT6
    generic map(
      INIT => X"AA2AAA2AFB3BFF3F"
    )
    port map (
      I0 => OVtpg_inst_pmode(2),
      I1 => OVtpg_inst_pmode(1),
      I2 => OVtpg_inst_pmode(0),
      I3 => N14,
      I4 => OVtpg_inst_Mmux_pixel_out_12_pixel_out_23_mux_50_OUT3166_296,
      I5 => OVtpg_inst_Mmux_pixel_out_12_pixel_out_23_mux_50_OUT3163_293,
      O => N130
    );
  OVtpg_inst_Active_glue_set : MUXF7
    port map (
      I0 => N136,
      I1 => N137,
      S => OVtpg_inst_n0315_inv1,
      O => OVtpg_inst_Active_glue_set_300
    );
  OVtpg_inst_Active_glue_set_F : LUT2
    generic map(
      INIT => X"B"
    )
    port map (
      I0 => OVtpg_inst_Active_235,
      I1 => locked_in,
      O => N136
    );
  OVtpg_inst_Active_glue_set_G : LUT6
    generic map(
      INIT => X"BBBBFBBBBBBBBBBB"
    )
    port map (
      I0 => OVtpg_inst_Active_235,
      I1 => locked_in,
      I2 => OVtpg_inst_Row_10_GND_7_o_equal_5_o_10_1_96,
      I3 => OVtpg_inst_Row(0),
      I4 => OVtpg_inst_Row(2),
      I5 => OVtpg_inst_Row(1),
      O => N137
    );
  OVtpg_inst_Row_10_PWR_7_o_div_45_o_0_14 : MUXF7
    port map (
      I0 => N138,
      I1 => N139,
      S => OVtpg_inst_Row_10_PWR_7_o_div_45_Madd_a_10_GND_9_o_add_19_OUT_10_0_lut_6_Q,
      O => OVtpg_inst_n0134(0)
    );
  OVtpg_inst_Row_10_PWR_7_o_div_45_o_0_14_F : LUT6
    generic map(
      INIT => X"AAA8A8A0A0808000"
    )
    port map (
      I0 => OVtpg_inst_Row_10_PWR_7_o_div_45_o_0_11,
      I1 => OVtpg_inst_Row_10_PWR_7_o_div_45_Madd_a_10_GND_9_o_add_19_OUT_10_0_lut_7_Q,
      I2 => OVtpg_inst_Row(4),
      I3 => OVtpg_inst_Row(2),
      I4 => OVtpg_inst_Row(3),
      I5 => OVtpg_inst_Row_10_PWR_7_o_div_45_n0441_8_Q,
      O => N138
    );
  OVtpg_inst_Row_10_PWR_7_o_div_45_o_0_14_G : LUT6
    generic map(
      INIT => X"2BA33FB7FFFFFFFF"
    )
    port map (
      I0 => OVtpg_inst_Row_10_PWR_7_o_div_45_Madd_a_10_GND_9_o_add_19_OUT_10_0_lut_7_Q,
      I1 => OVtpg_inst_Row(4),
      I2 => OVtpg_inst_Row_10_PWR_7_o_div_45_n0441_8_Q,
      I3 => OVtpg_inst_Row_10_PWR_7_o_div_45_o_0_12,
      I4 => OVtpg_inst_Row(3),
      I5 => OVtpg_inst_Row_10_PWR_7_o_div_45_o_0_11,
      O => N139
    );
  OVtpg_inst_Mmux_pixel_out_12_pixel_out_23_mux_50_OUT31611_SW0 : MUXF7
    port map (
      I0 => N140,
      I1 => N141,
      S => OVtpg_inst_Row_10_PWR_7_o_div_45_o_0_11,
      O => N22
    );
  OVtpg_inst_Mmux_pixel_out_12_pixel_out_23_mux_50_OUT31611_SW0_G : LUT6
    generic map(
      INIT => X"4555155523111555"
    )
    port map (
      I0 => OVtpg_inst_Row_10_PWR_7_o_div_45_Madd_a_10_GND_9_o_add_19_OUT_10_0_lut_7_Q,
      I1 => OVtpg_inst_Row_10_PWR_7_o_div_45_n0441_8_Q,
      I2 => OVtpg_inst_Row(3),
      I3 => OVtpg_inst_Row_10_PWR_7_o_div_45_Madd_a_10_GND_9_o_add_19_OUT_10_0_lut_6_Q,
      I4 => OVtpg_inst_Row(4),
      I5 => OVtpg_inst_Row_10_PWR_7_o_div_45_o_0_12,
      O => N141
    );
  OVtpg_inst_Vsynci_glue_set_G : LUT6
    generic map(
      INIT => X"AA8AAAAAAABAAAAA"
    )
    port map (
      I0 => OVtpg_inst_Vsynci_237,
      I1 => OVtpg_inst_Row(4),
      I2 => OVtpg_inst_Row_10_GND_7_o_equal_8_o_10_1,
      I3 => OVtpg_inst_Row(2),
      I4 => OVtpg_inst_Row(5),
      I5 => OVtpg_inst_Row(1),
      O => N143
    );
  OVtpg_inst_Mcount_Col_lut_0_INV_0 : INV
    port map (
      I => OVtpg_inst_Col(0),
      O => OVtpg_inst_Mcount_Col_lut(0)
    );
  OVtpg_inst_Mcount_Row_lut_0_INV_0 : INV
    port map (
      I => OVtpg_inst_Row(0),
      O => OVtpg_inst_Mcount_Row_lut(0)
    );
  OVtpg_inst_Mcount_addr_lut_0_INV_0 : INV
    port map (
      I => NlwRenamedSig_OI_OVtpg_inst_addr(0),
      O => OVtpg_inst_Mcount_addr_lut(0)
    );
  MRST1_INV_0 : INV
    port map (
      I => locked_in,
      O => MRST
    );
  OVtpg_inst_PCLK1_INV_0 : INV
    port map (
      I => OVtpg_inst_ClkDiv(0),
      O => OVtpg_inst_PCLK
    );
  SIF_inst_oddpix_INV_358_o1_INV_0 : INV
    port map (
      I => SIF_inst_oddpix_252,
      O => SIF_inst_oddpix_INV_358_o
    );
  SIF_inst_VS_in_INV_360_o1_INV_0 : INV
    port map (
      I => OVtpg_inst_VSYNC_60,
      O => SIF_inst_VS_in_INV_360_o
    );
  Vsync_inv1_INV_0 : INV
    port map (
      I => NlwRenamedSig_OI_SIF_inst_Vsync,
      O => vid_vsync
    );
  Hsync_inv1_INV_0 : INV
    port map (
      I => NlwRenamedSig_OI_SIF_inst_Hsync,
      O => vid_hsync
    );
  OVtpg_inst_Mmux_pixel_out_12_pixel_out_23_mux_50_OUT31611_SW0_F_INV_0 : INV
    port map (
      I => OVtpg_inst_Row_10_PWR_7_o_div_45_Madd_a_10_GND_9_o_add_19_OUT_10_0_lut_7_Q,
      O => N140
    );
  OVtpg_inst_Vsynci_glue_set1 : LUT3
    generic map(
      INIT => X"E4"
    )
    port map (
      I0 => OVtpg_inst_n0315_inv1,
      I1 => OVtpg_inst_Vsynci_237,
      I2 => N143,
      O => OVtpg_inst_Vsynci_glue_set
    );

end Structure;
